VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 1760.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 42.560 2800.000 43.120 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1280.160 4.000 1280.720 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1061.760 4.000 1062.320 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 843.360 4.000 843.920 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 624.960 4.000 625.520 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 406.560 4.000 407.120 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 188.160 4.000 188.720 ;
    END
  END io_in[15]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 260.960 2800.000 261.520 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 479.360 2800.000 479.920 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 697.760 2800.000 698.320 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 916.160 2800.000 916.720 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1134.560 2800.000 1135.120 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1352.960 2800.000 1353.520 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1571.360 2800.000 1571.920 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1716.960 4.000 1717.520 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1498.560 4.000 1499.120 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 188.160 2800.000 188.720 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1134.560 4.000 1135.120 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 916.160 4.000 916.720 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 697.760 4.000 698.320 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 479.360 4.000 479.920 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 260.960 4.000 261.520 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 42.560 4.000 43.120 ;
    END
  END io_oeb[15]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 406.560 2800.000 407.120 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 624.960 2800.000 625.520 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 843.360 2800.000 843.920 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1061.760 2800.000 1062.320 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1280.160 2800.000 1280.720 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1498.560 2800.000 1499.120 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1716.960 2800.000 1717.520 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1571.360 4.000 1571.920 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1352.960 4.000 1353.520 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 115.360 2800.000 115.920 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1207.360 4.000 1207.920 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 988.960 4.000 989.520 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 770.560 4.000 771.120 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 552.160 4.000 552.720 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 333.760 4.000 334.320 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 115.360 4.000 115.920 ;
    END
  END io_out[15]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 333.760 2800.000 334.320 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 552.160 2800.000 552.720 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 770.560 2800.000 771.120 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 988.960 2800.000 989.520 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1207.360 2800.000 1207.920 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1425.760 2800.000 1426.320 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2796.000 1644.160 2800.000 1644.720 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1644.160 4.000 1644.720 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1425.760 4.000 1426.320 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2765.840 0.000 2766.400 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2771.440 0.000 2772.000 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2777.040 0.000 2777.600 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 615.440 0.000 616.000 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2295.440 0.000 2296.000 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2312.240 0.000 2312.800 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2329.040 0.000 2329.600 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2345.840 0.000 2346.400 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2362.640 0.000 2363.200 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2379.440 0.000 2380.000 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2396.240 0.000 2396.800 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2413.040 0.000 2413.600 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2429.840 0.000 2430.400 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2446.640 0.000 2447.200 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 783.440 0.000 784.000 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2463.440 0.000 2464.000 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2480.240 0.000 2480.800 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2497.040 0.000 2497.600 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2513.840 0.000 2514.400 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2530.640 0.000 2531.200 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2547.440 0.000 2548.000 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2564.240 0.000 2564.800 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2581.040 0.000 2581.600 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2597.840 0.000 2598.400 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2614.640 0.000 2615.200 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 800.240 0.000 800.800 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2631.440 0.000 2632.000 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2648.240 0.000 2648.800 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2665.040 0.000 2665.600 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2681.840 0.000 2682.400 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2698.640 0.000 2699.200 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2715.440 0.000 2716.000 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2732.240 0.000 2732.800 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2749.040 0.000 2749.600 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 817.040 0.000 817.600 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 833.840 0.000 834.400 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 850.640 0.000 851.200 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 867.440 0.000 868.000 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 884.240 0.000 884.800 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 901.040 0.000 901.600 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 917.840 0.000 918.400 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 934.640 0.000 935.200 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 632.240 0.000 632.800 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 951.440 0.000 952.000 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 968.240 0.000 968.800 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 985.040 0.000 985.600 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1001.840 0.000 1002.400 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1018.640 0.000 1019.200 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1035.440 0.000 1036.000 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1052.240 0.000 1052.800 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1069.040 0.000 1069.600 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1085.840 0.000 1086.400 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1102.640 0.000 1103.200 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 649.040 0.000 649.600 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1119.440 0.000 1120.000 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1136.240 0.000 1136.800 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1153.040 0.000 1153.600 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1169.840 0.000 1170.400 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1186.640 0.000 1187.200 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1203.440 0.000 1204.000 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1220.240 0.000 1220.800 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1237.040 0.000 1237.600 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1253.840 0.000 1254.400 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1270.640 0.000 1271.200 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 665.840 0.000 666.400 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1287.440 0.000 1288.000 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1304.240 0.000 1304.800 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1321.040 0.000 1321.600 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1337.840 0.000 1338.400 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1354.640 0.000 1355.200 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1371.440 0.000 1372.000 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1388.240 0.000 1388.800 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1405.040 0.000 1405.600 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1421.840 0.000 1422.400 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1438.640 0.000 1439.200 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 682.640 0.000 683.200 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1455.440 0.000 1456.000 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1472.240 0.000 1472.800 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1489.040 0.000 1489.600 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1505.840 0.000 1506.400 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1522.640 0.000 1523.200 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1539.440 0.000 1540.000 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1556.240 0.000 1556.800 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1573.040 0.000 1573.600 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1589.840 0.000 1590.400 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1606.640 0.000 1607.200 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 699.440 0.000 700.000 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1623.440 0.000 1624.000 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1640.240 0.000 1640.800 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1657.040 0.000 1657.600 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1673.840 0.000 1674.400 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1690.640 0.000 1691.200 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1707.440 0.000 1708.000 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1724.240 0.000 1724.800 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1741.040 0.000 1741.600 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1757.840 0.000 1758.400 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1774.640 0.000 1775.200 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 716.240 0.000 716.800 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1791.440 0.000 1792.000 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1808.240 0.000 1808.800 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1825.040 0.000 1825.600 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1841.840 0.000 1842.400 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1858.640 0.000 1859.200 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1875.440 0.000 1876.000 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1892.240 0.000 1892.800 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1909.040 0.000 1909.600 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1925.840 0.000 1926.400 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1942.640 0.000 1943.200 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 733.040 0.000 733.600 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1959.440 0.000 1960.000 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1976.240 0.000 1976.800 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1993.040 0.000 1993.600 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2009.840 0.000 2010.400 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2026.640 0.000 2027.200 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2043.440 0.000 2044.000 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2060.240 0.000 2060.800 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2077.040 0.000 2077.600 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2093.840 0.000 2094.400 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2110.640 0.000 2111.200 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 749.840 0.000 750.400 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2127.440 0.000 2128.000 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2144.240 0.000 2144.800 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2161.040 0.000 2161.600 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2177.840 0.000 2178.400 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2194.640 0.000 2195.200 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2211.440 0.000 2212.000 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2228.240 0.000 2228.800 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2245.040 0.000 2245.600 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2261.840 0.000 2262.400 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2278.640 0.000 2279.200 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 766.640 0.000 767.200 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 621.040 0.000 621.600 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2301.040 0.000 2301.600 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2317.840 0.000 2318.400 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2334.640 0.000 2335.200 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2351.440 0.000 2352.000 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2368.240 0.000 2368.800 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2385.040 0.000 2385.600 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2401.840 0.000 2402.400 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2418.640 0.000 2419.200 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2435.440 0.000 2436.000 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2452.240 0.000 2452.800 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 789.040 0.000 789.600 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2469.040 0.000 2469.600 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2485.840 0.000 2486.400 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2502.640 0.000 2503.200 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2519.440 0.000 2520.000 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2536.240 0.000 2536.800 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2553.040 0.000 2553.600 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2569.840 0.000 2570.400 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2586.640 0.000 2587.200 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2603.440 0.000 2604.000 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2620.240 0.000 2620.800 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 805.840 0.000 806.400 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2637.040 0.000 2637.600 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2653.840 0.000 2654.400 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2670.640 0.000 2671.200 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2687.440 0.000 2688.000 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2704.240 0.000 2704.800 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2721.040 0.000 2721.600 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2737.840 0.000 2738.400 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2754.640 0.000 2755.200 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 822.640 0.000 823.200 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 839.440 0.000 840.000 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 856.240 0.000 856.800 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 873.040 0.000 873.600 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 889.840 0.000 890.400 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 906.640 0.000 907.200 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 923.440 0.000 924.000 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 940.240 0.000 940.800 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 637.840 0.000 638.400 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 957.040 0.000 957.600 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 973.840 0.000 974.400 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 990.640 0.000 991.200 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1007.440 0.000 1008.000 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1024.240 0.000 1024.800 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1041.040 0.000 1041.600 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1057.840 0.000 1058.400 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1074.640 0.000 1075.200 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1091.440 0.000 1092.000 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1108.240 0.000 1108.800 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 654.640 0.000 655.200 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1125.040 0.000 1125.600 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1141.840 0.000 1142.400 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1158.640 0.000 1159.200 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1175.440 0.000 1176.000 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1192.240 0.000 1192.800 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1209.040 0.000 1209.600 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1225.840 0.000 1226.400 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1242.640 0.000 1243.200 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1259.440 0.000 1260.000 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1276.240 0.000 1276.800 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 671.440 0.000 672.000 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1293.040 0.000 1293.600 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1309.840 0.000 1310.400 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1326.640 0.000 1327.200 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1343.440 0.000 1344.000 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1360.240 0.000 1360.800 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1377.040 0.000 1377.600 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1393.840 0.000 1394.400 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1410.640 0.000 1411.200 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1427.440 0.000 1428.000 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1444.240 0.000 1444.800 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 688.240 0.000 688.800 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1461.040 0.000 1461.600 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1477.840 0.000 1478.400 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1494.640 0.000 1495.200 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1511.440 0.000 1512.000 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1528.240 0.000 1528.800 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1545.040 0.000 1545.600 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1561.840 0.000 1562.400 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1578.640 0.000 1579.200 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1595.440 0.000 1596.000 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1612.240 0.000 1612.800 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 705.040 0.000 705.600 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1629.040 0.000 1629.600 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1645.840 0.000 1646.400 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1662.640 0.000 1663.200 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1679.440 0.000 1680.000 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1696.240 0.000 1696.800 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1713.040 0.000 1713.600 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1729.840 0.000 1730.400 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1746.640 0.000 1747.200 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1763.440 0.000 1764.000 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1780.240 0.000 1780.800 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 721.840 0.000 722.400 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1797.040 0.000 1797.600 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1813.840 0.000 1814.400 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1830.640 0.000 1831.200 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1847.440 0.000 1848.000 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1864.240 0.000 1864.800 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1881.040 0.000 1881.600 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1897.840 0.000 1898.400 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1914.640 0.000 1915.200 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1931.440 0.000 1932.000 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1948.240 0.000 1948.800 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 738.640 0.000 739.200 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1965.040 0.000 1965.600 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1981.840 0.000 1982.400 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1998.640 0.000 1999.200 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2015.440 0.000 2016.000 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2032.240 0.000 2032.800 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2049.040 0.000 2049.600 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2065.840 0.000 2066.400 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2082.640 0.000 2083.200 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2099.440 0.000 2100.000 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2116.240 0.000 2116.800 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 755.440 0.000 756.000 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2133.040 0.000 2133.600 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2149.840 0.000 2150.400 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2166.640 0.000 2167.200 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2183.440 0.000 2184.000 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2200.240 0.000 2200.800 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2217.040 0.000 2217.600 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2233.840 0.000 2234.400 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2250.640 0.000 2251.200 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2267.440 0.000 2268.000 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2284.240 0.000 2284.800 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 772.240 0.000 772.800 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 626.640 0.000 627.200 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2306.640 0.000 2307.200 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2323.440 0.000 2324.000 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2340.240 0.000 2340.800 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2357.040 0.000 2357.600 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2373.840 0.000 2374.400 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2390.640 0.000 2391.200 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2407.440 0.000 2408.000 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2424.240 0.000 2424.800 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2441.040 0.000 2441.600 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2457.840 0.000 2458.400 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 794.640 0.000 795.200 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2474.640 0.000 2475.200 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2491.440 0.000 2492.000 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2508.240 0.000 2508.800 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2525.040 0.000 2525.600 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2541.840 0.000 2542.400 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2558.640 0.000 2559.200 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2575.440 0.000 2576.000 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2592.240 0.000 2592.800 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2609.040 0.000 2609.600 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2625.840 0.000 2626.400 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 811.440 0.000 812.000 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2642.640 0.000 2643.200 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2659.440 0.000 2660.000 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2676.240 0.000 2676.800 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2693.040 0.000 2693.600 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2709.840 0.000 2710.400 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2726.640 0.000 2727.200 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2743.440 0.000 2744.000 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2760.240 0.000 2760.800 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 828.240 0.000 828.800 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 845.040 0.000 845.600 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 861.840 0.000 862.400 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 878.640 0.000 879.200 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 895.440 0.000 896.000 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 912.240 0.000 912.800 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 929.040 0.000 929.600 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 945.840 0.000 946.400 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 643.440 0.000 644.000 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 962.640 0.000 963.200 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 979.440 0.000 980.000 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 996.240 0.000 996.800 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1013.040 0.000 1013.600 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1029.840 0.000 1030.400 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1046.640 0.000 1047.200 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1063.440 0.000 1064.000 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1080.240 0.000 1080.800 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1097.040 0.000 1097.600 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1113.840 0.000 1114.400 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 660.240 0.000 660.800 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1130.640 0.000 1131.200 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1147.440 0.000 1148.000 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1164.240 0.000 1164.800 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1181.040 0.000 1181.600 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1197.840 0.000 1198.400 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1214.640 0.000 1215.200 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1231.440 0.000 1232.000 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1248.240 0.000 1248.800 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1265.040 0.000 1265.600 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1281.840 0.000 1282.400 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 677.040 0.000 677.600 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1298.640 0.000 1299.200 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1315.440 0.000 1316.000 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1332.240 0.000 1332.800 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1349.040 0.000 1349.600 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1365.840 0.000 1366.400 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1382.640 0.000 1383.200 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1399.440 0.000 1400.000 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1416.240 0.000 1416.800 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1433.040 0.000 1433.600 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1449.840 0.000 1450.400 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 693.840 0.000 694.400 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1466.640 0.000 1467.200 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1483.440 0.000 1484.000 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1500.240 0.000 1500.800 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1517.040 0.000 1517.600 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1533.840 0.000 1534.400 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1550.640 0.000 1551.200 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1567.440 0.000 1568.000 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1584.240 0.000 1584.800 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1601.040 0.000 1601.600 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1617.840 0.000 1618.400 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 710.640 0.000 711.200 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1634.640 0.000 1635.200 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1651.440 0.000 1652.000 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1668.240 0.000 1668.800 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1685.040 0.000 1685.600 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1701.840 0.000 1702.400 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1718.640 0.000 1719.200 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1735.440 0.000 1736.000 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1752.240 0.000 1752.800 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1769.040 0.000 1769.600 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1785.840 0.000 1786.400 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 727.440 0.000 728.000 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1802.640 0.000 1803.200 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1819.440 0.000 1820.000 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1836.240 0.000 1836.800 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1853.040 0.000 1853.600 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1869.840 0.000 1870.400 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1886.640 0.000 1887.200 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1903.440 0.000 1904.000 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1920.240 0.000 1920.800 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1937.040 0.000 1937.600 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1953.840 0.000 1954.400 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 744.240 0.000 744.800 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1970.640 0.000 1971.200 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1987.440 0.000 1988.000 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2004.240 0.000 2004.800 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2021.040 0.000 2021.600 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2037.840 0.000 2038.400 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2054.640 0.000 2055.200 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2071.440 0.000 2072.000 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2088.240 0.000 2088.800 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2105.040 0.000 2105.600 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2121.840 0.000 2122.400 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 761.040 0.000 761.600 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2138.640 0.000 2139.200 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2155.440 0.000 2156.000 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2172.240 0.000 2172.800 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2189.040 0.000 2189.600 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2205.840 0.000 2206.400 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2222.640 0.000 2223.200 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2239.440 0.000 2240.000 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2256.240 0.000 2256.800 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2273.040 0.000 2273.600 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2289.840 0.000 2290.400 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 777.840 0.000 778.400 4.000 ;
    END
  END la_oenb[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 15.380 1406.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1558.240 15.380 1559.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1711.840 15.380 1713.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1865.440 15.380 1867.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2019.040 15.380 2020.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2172.640 15.380 2174.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2326.240 15.380 2327.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2479.840 15.380 2481.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2633.440 15.380 2635.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2787.040 15.380 2788.640 1740.780 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.840 15.380 1329.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1481.440 15.380 1483.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.040 15.380 1636.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1788.640 15.380 1790.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1942.240 15.380 1943.840 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2095.840 15.380 2097.440 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2249.440 15.380 2251.040 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2403.040 15.380 2404.640 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2556.640 15.380 2558.240 1740.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2710.240 15.380 2711.840 1740.780 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 21.840 0.000 22.400 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 27.440 0.000 28.000 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.040 0.000 33.600 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 55.440 0.000 56.000 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 245.840 0.000 246.400 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.640 0.000 263.200 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 279.440 0.000 280.000 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 296.240 0.000 296.800 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 313.040 0.000 313.600 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.840 0.000 330.400 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 346.640 0.000 347.200 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 363.440 0.000 364.000 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 380.240 0.000 380.800 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 397.040 0.000 397.600 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.840 0.000 78.400 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 413.840 0.000 414.400 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 430.640 0.000 431.200 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 447.440 0.000 448.000 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 464.240 0.000 464.800 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 481.040 0.000 481.600 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.840 0.000 498.400 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 514.640 0.000 515.200 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 531.440 0.000 532.000 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 548.240 0.000 548.800 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 565.040 0.000 565.600 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.240 0.000 100.800 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 581.840 0.000 582.400 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 598.640 0.000 599.200 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 122.640 0.000 123.200 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 145.040 0.000 145.600 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.840 0.000 162.400 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 178.640 0.000 179.200 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 195.440 0.000 196.000 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 212.240 0.000 212.800 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 229.040 0.000 229.600 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 38.640 0.000 39.200 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 61.040 0.000 61.600 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 251.440 0.000 252.000 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.240 0.000 268.800 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 285.040 0.000 285.600 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 301.840 0.000 302.400 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 318.640 0.000 319.200 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 335.440 0.000 336.000 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 352.240 0.000 352.800 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 369.040 0.000 369.600 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 385.840 0.000 386.400 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 402.640 0.000 403.200 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 83.440 0.000 84.000 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 419.440 0.000 420.000 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 436.240 0.000 436.800 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 453.040 0.000 453.600 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 469.840 0.000 470.400 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 486.640 0.000 487.200 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 503.440 0.000 504.000 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 520.240 0.000 520.800 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 537.040 0.000 537.600 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 553.840 0.000 554.400 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 570.640 0.000 571.200 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 105.840 0.000 106.400 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 587.440 0.000 588.000 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 604.240 0.000 604.800 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 128.240 0.000 128.800 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 150.640 0.000 151.200 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 167.440 0.000 168.000 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.240 0.000 184.800 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.040 0.000 201.600 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 217.840 0.000 218.400 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.640 0.000 235.200 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.640 0.000 67.200 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 257.040 0.000 257.600 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 273.840 0.000 274.400 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 290.640 0.000 291.200 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 307.440 0.000 308.000 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 324.240 0.000 324.800 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 341.040 0.000 341.600 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 357.840 0.000 358.400 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 374.640 0.000 375.200 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 391.440 0.000 392.000 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 408.240 0.000 408.800 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 89.040 0.000 89.600 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 425.040 0.000 425.600 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 441.840 0.000 442.400 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 458.640 0.000 459.200 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 475.440 0.000 476.000 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 492.240 0.000 492.800 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 509.040 0.000 509.600 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 525.840 0.000 526.400 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 542.640 0.000 543.200 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 559.440 0.000 560.000 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 576.240 0.000 576.800 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 111.440 0.000 112.000 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 593.040 0.000 593.600 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 609.840 0.000 610.400 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 133.840 0.000 134.400 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 156.240 0.000 156.800 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 173.040 0.000 173.600 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 189.840 0.000 190.400 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 206.640 0.000 207.200 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 223.440 0.000 224.000 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 240.240 0.000 240.800 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 72.240 0.000 72.800 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.640 0.000 95.200 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.040 0.000 117.600 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 139.440 0.000 140.000 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 44.240 0.000 44.800 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 49.840 0.000 50.400 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 8.550 2793.280 1740.780 ;
      LAYER Metal2 ;
        RECT 4.620 4.300 2792.580 1740.670 ;
        RECT 4.620 2.890 21.540 4.300 ;
        RECT 22.700 2.890 27.140 4.300 ;
        RECT 28.300 2.890 32.740 4.300 ;
        RECT 33.900 2.890 38.340 4.300 ;
        RECT 39.500 2.890 43.940 4.300 ;
        RECT 45.100 2.890 49.540 4.300 ;
        RECT 50.700 2.890 55.140 4.300 ;
        RECT 56.300 2.890 60.740 4.300 ;
        RECT 61.900 2.890 66.340 4.300 ;
        RECT 67.500 2.890 71.940 4.300 ;
        RECT 73.100 2.890 77.540 4.300 ;
        RECT 78.700 2.890 83.140 4.300 ;
        RECT 84.300 2.890 88.740 4.300 ;
        RECT 89.900 2.890 94.340 4.300 ;
        RECT 95.500 2.890 99.940 4.300 ;
        RECT 101.100 2.890 105.540 4.300 ;
        RECT 106.700 2.890 111.140 4.300 ;
        RECT 112.300 2.890 116.740 4.300 ;
        RECT 117.900 2.890 122.340 4.300 ;
        RECT 123.500 2.890 127.940 4.300 ;
        RECT 129.100 2.890 133.540 4.300 ;
        RECT 134.700 2.890 139.140 4.300 ;
        RECT 140.300 2.890 144.740 4.300 ;
        RECT 145.900 2.890 150.340 4.300 ;
        RECT 151.500 2.890 155.940 4.300 ;
        RECT 157.100 2.890 161.540 4.300 ;
        RECT 162.700 2.890 167.140 4.300 ;
        RECT 168.300 2.890 172.740 4.300 ;
        RECT 173.900 2.890 178.340 4.300 ;
        RECT 179.500 2.890 183.940 4.300 ;
        RECT 185.100 2.890 189.540 4.300 ;
        RECT 190.700 2.890 195.140 4.300 ;
        RECT 196.300 2.890 200.740 4.300 ;
        RECT 201.900 2.890 206.340 4.300 ;
        RECT 207.500 2.890 211.940 4.300 ;
        RECT 213.100 2.890 217.540 4.300 ;
        RECT 218.700 2.890 223.140 4.300 ;
        RECT 224.300 2.890 228.740 4.300 ;
        RECT 229.900 2.890 234.340 4.300 ;
        RECT 235.500 2.890 239.940 4.300 ;
        RECT 241.100 2.890 245.540 4.300 ;
        RECT 246.700 2.890 251.140 4.300 ;
        RECT 252.300 2.890 256.740 4.300 ;
        RECT 257.900 2.890 262.340 4.300 ;
        RECT 263.500 2.890 267.940 4.300 ;
        RECT 269.100 2.890 273.540 4.300 ;
        RECT 274.700 2.890 279.140 4.300 ;
        RECT 280.300 2.890 284.740 4.300 ;
        RECT 285.900 2.890 290.340 4.300 ;
        RECT 291.500 2.890 295.940 4.300 ;
        RECT 297.100 2.890 301.540 4.300 ;
        RECT 302.700 2.890 307.140 4.300 ;
        RECT 308.300 2.890 312.740 4.300 ;
        RECT 313.900 2.890 318.340 4.300 ;
        RECT 319.500 2.890 323.940 4.300 ;
        RECT 325.100 2.890 329.540 4.300 ;
        RECT 330.700 2.890 335.140 4.300 ;
        RECT 336.300 2.890 340.740 4.300 ;
        RECT 341.900 2.890 346.340 4.300 ;
        RECT 347.500 2.890 351.940 4.300 ;
        RECT 353.100 2.890 357.540 4.300 ;
        RECT 358.700 2.890 363.140 4.300 ;
        RECT 364.300 2.890 368.740 4.300 ;
        RECT 369.900 2.890 374.340 4.300 ;
        RECT 375.500 2.890 379.940 4.300 ;
        RECT 381.100 2.890 385.540 4.300 ;
        RECT 386.700 2.890 391.140 4.300 ;
        RECT 392.300 2.890 396.740 4.300 ;
        RECT 397.900 2.890 402.340 4.300 ;
        RECT 403.500 2.890 407.940 4.300 ;
        RECT 409.100 2.890 413.540 4.300 ;
        RECT 414.700 2.890 419.140 4.300 ;
        RECT 420.300 2.890 424.740 4.300 ;
        RECT 425.900 2.890 430.340 4.300 ;
        RECT 431.500 2.890 435.940 4.300 ;
        RECT 437.100 2.890 441.540 4.300 ;
        RECT 442.700 2.890 447.140 4.300 ;
        RECT 448.300 2.890 452.740 4.300 ;
        RECT 453.900 2.890 458.340 4.300 ;
        RECT 459.500 2.890 463.940 4.300 ;
        RECT 465.100 2.890 469.540 4.300 ;
        RECT 470.700 2.890 475.140 4.300 ;
        RECT 476.300 2.890 480.740 4.300 ;
        RECT 481.900 2.890 486.340 4.300 ;
        RECT 487.500 2.890 491.940 4.300 ;
        RECT 493.100 2.890 497.540 4.300 ;
        RECT 498.700 2.890 503.140 4.300 ;
        RECT 504.300 2.890 508.740 4.300 ;
        RECT 509.900 2.890 514.340 4.300 ;
        RECT 515.500 2.890 519.940 4.300 ;
        RECT 521.100 2.890 525.540 4.300 ;
        RECT 526.700 2.890 531.140 4.300 ;
        RECT 532.300 2.890 536.740 4.300 ;
        RECT 537.900 2.890 542.340 4.300 ;
        RECT 543.500 2.890 547.940 4.300 ;
        RECT 549.100 2.890 553.540 4.300 ;
        RECT 554.700 2.890 559.140 4.300 ;
        RECT 560.300 2.890 564.740 4.300 ;
        RECT 565.900 2.890 570.340 4.300 ;
        RECT 571.500 2.890 575.940 4.300 ;
        RECT 577.100 2.890 581.540 4.300 ;
        RECT 582.700 2.890 587.140 4.300 ;
        RECT 588.300 2.890 592.740 4.300 ;
        RECT 593.900 2.890 598.340 4.300 ;
        RECT 599.500 2.890 603.940 4.300 ;
        RECT 605.100 2.890 609.540 4.300 ;
        RECT 610.700 2.890 615.140 4.300 ;
        RECT 616.300 2.890 620.740 4.300 ;
        RECT 621.900 2.890 626.340 4.300 ;
        RECT 627.500 2.890 631.940 4.300 ;
        RECT 633.100 2.890 637.540 4.300 ;
        RECT 638.700 2.890 643.140 4.300 ;
        RECT 644.300 2.890 648.740 4.300 ;
        RECT 649.900 2.890 654.340 4.300 ;
        RECT 655.500 2.890 659.940 4.300 ;
        RECT 661.100 2.890 665.540 4.300 ;
        RECT 666.700 2.890 671.140 4.300 ;
        RECT 672.300 2.890 676.740 4.300 ;
        RECT 677.900 2.890 682.340 4.300 ;
        RECT 683.500 2.890 687.940 4.300 ;
        RECT 689.100 2.890 693.540 4.300 ;
        RECT 694.700 2.890 699.140 4.300 ;
        RECT 700.300 2.890 704.740 4.300 ;
        RECT 705.900 2.890 710.340 4.300 ;
        RECT 711.500 2.890 715.940 4.300 ;
        RECT 717.100 2.890 721.540 4.300 ;
        RECT 722.700 2.890 727.140 4.300 ;
        RECT 728.300 2.890 732.740 4.300 ;
        RECT 733.900 2.890 738.340 4.300 ;
        RECT 739.500 2.890 743.940 4.300 ;
        RECT 745.100 2.890 749.540 4.300 ;
        RECT 750.700 2.890 755.140 4.300 ;
        RECT 756.300 2.890 760.740 4.300 ;
        RECT 761.900 2.890 766.340 4.300 ;
        RECT 767.500 2.890 771.940 4.300 ;
        RECT 773.100 2.890 777.540 4.300 ;
        RECT 778.700 2.890 783.140 4.300 ;
        RECT 784.300 2.890 788.740 4.300 ;
        RECT 789.900 2.890 794.340 4.300 ;
        RECT 795.500 2.890 799.940 4.300 ;
        RECT 801.100 2.890 805.540 4.300 ;
        RECT 806.700 2.890 811.140 4.300 ;
        RECT 812.300 2.890 816.740 4.300 ;
        RECT 817.900 2.890 822.340 4.300 ;
        RECT 823.500 2.890 827.940 4.300 ;
        RECT 829.100 2.890 833.540 4.300 ;
        RECT 834.700 2.890 839.140 4.300 ;
        RECT 840.300 2.890 844.740 4.300 ;
        RECT 845.900 2.890 850.340 4.300 ;
        RECT 851.500 2.890 855.940 4.300 ;
        RECT 857.100 2.890 861.540 4.300 ;
        RECT 862.700 2.890 867.140 4.300 ;
        RECT 868.300 2.890 872.740 4.300 ;
        RECT 873.900 2.890 878.340 4.300 ;
        RECT 879.500 2.890 883.940 4.300 ;
        RECT 885.100 2.890 889.540 4.300 ;
        RECT 890.700 2.890 895.140 4.300 ;
        RECT 896.300 2.890 900.740 4.300 ;
        RECT 901.900 2.890 906.340 4.300 ;
        RECT 907.500 2.890 911.940 4.300 ;
        RECT 913.100 2.890 917.540 4.300 ;
        RECT 918.700 2.890 923.140 4.300 ;
        RECT 924.300 2.890 928.740 4.300 ;
        RECT 929.900 2.890 934.340 4.300 ;
        RECT 935.500 2.890 939.940 4.300 ;
        RECT 941.100 2.890 945.540 4.300 ;
        RECT 946.700 2.890 951.140 4.300 ;
        RECT 952.300 2.890 956.740 4.300 ;
        RECT 957.900 2.890 962.340 4.300 ;
        RECT 963.500 2.890 967.940 4.300 ;
        RECT 969.100 2.890 973.540 4.300 ;
        RECT 974.700 2.890 979.140 4.300 ;
        RECT 980.300 2.890 984.740 4.300 ;
        RECT 985.900 2.890 990.340 4.300 ;
        RECT 991.500 2.890 995.940 4.300 ;
        RECT 997.100 2.890 1001.540 4.300 ;
        RECT 1002.700 2.890 1007.140 4.300 ;
        RECT 1008.300 2.890 1012.740 4.300 ;
        RECT 1013.900 2.890 1018.340 4.300 ;
        RECT 1019.500 2.890 1023.940 4.300 ;
        RECT 1025.100 2.890 1029.540 4.300 ;
        RECT 1030.700 2.890 1035.140 4.300 ;
        RECT 1036.300 2.890 1040.740 4.300 ;
        RECT 1041.900 2.890 1046.340 4.300 ;
        RECT 1047.500 2.890 1051.940 4.300 ;
        RECT 1053.100 2.890 1057.540 4.300 ;
        RECT 1058.700 2.890 1063.140 4.300 ;
        RECT 1064.300 2.890 1068.740 4.300 ;
        RECT 1069.900 2.890 1074.340 4.300 ;
        RECT 1075.500 2.890 1079.940 4.300 ;
        RECT 1081.100 2.890 1085.540 4.300 ;
        RECT 1086.700 2.890 1091.140 4.300 ;
        RECT 1092.300 2.890 1096.740 4.300 ;
        RECT 1097.900 2.890 1102.340 4.300 ;
        RECT 1103.500 2.890 1107.940 4.300 ;
        RECT 1109.100 2.890 1113.540 4.300 ;
        RECT 1114.700 2.890 1119.140 4.300 ;
        RECT 1120.300 2.890 1124.740 4.300 ;
        RECT 1125.900 2.890 1130.340 4.300 ;
        RECT 1131.500 2.890 1135.940 4.300 ;
        RECT 1137.100 2.890 1141.540 4.300 ;
        RECT 1142.700 2.890 1147.140 4.300 ;
        RECT 1148.300 2.890 1152.740 4.300 ;
        RECT 1153.900 2.890 1158.340 4.300 ;
        RECT 1159.500 2.890 1163.940 4.300 ;
        RECT 1165.100 2.890 1169.540 4.300 ;
        RECT 1170.700 2.890 1175.140 4.300 ;
        RECT 1176.300 2.890 1180.740 4.300 ;
        RECT 1181.900 2.890 1186.340 4.300 ;
        RECT 1187.500 2.890 1191.940 4.300 ;
        RECT 1193.100 2.890 1197.540 4.300 ;
        RECT 1198.700 2.890 1203.140 4.300 ;
        RECT 1204.300 2.890 1208.740 4.300 ;
        RECT 1209.900 2.890 1214.340 4.300 ;
        RECT 1215.500 2.890 1219.940 4.300 ;
        RECT 1221.100 2.890 1225.540 4.300 ;
        RECT 1226.700 2.890 1231.140 4.300 ;
        RECT 1232.300 2.890 1236.740 4.300 ;
        RECT 1237.900 2.890 1242.340 4.300 ;
        RECT 1243.500 2.890 1247.940 4.300 ;
        RECT 1249.100 2.890 1253.540 4.300 ;
        RECT 1254.700 2.890 1259.140 4.300 ;
        RECT 1260.300 2.890 1264.740 4.300 ;
        RECT 1265.900 2.890 1270.340 4.300 ;
        RECT 1271.500 2.890 1275.940 4.300 ;
        RECT 1277.100 2.890 1281.540 4.300 ;
        RECT 1282.700 2.890 1287.140 4.300 ;
        RECT 1288.300 2.890 1292.740 4.300 ;
        RECT 1293.900 2.890 1298.340 4.300 ;
        RECT 1299.500 2.890 1303.940 4.300 ;
        RECT 1305.100 2.890 1309.540 4.300 ;
        RECT 1310.700 2.890 1315.140 4.300 ;
        RECT 1316.300 2.890 1320.740 4.300 ;
        RECT 1321.900 2.890 1326.340 4.300 ;
        RECT 1327.500 2.890 1331.940 4.300 ;
        RECT 1333.100 2.890 1337.540 4.300 ;
        RECT 1338.700 2.890 1343.140 4.300 ;
        RECT 1344.300 2.890 1348.740 4.300 ;
        RECT 1349.900 2.890 1354.340 4.300 ;
        RECT 1355.500 2.890 1359.940 4.300 ;
        RECT 1361.100 2.890 1365.540 4.300 ;
        RECT 1366.700 2.890 1371.140 4.300 ;
        RECT 1372.300 2.890 1376.740 4.300 ;
        RECT 1377.900 2.890 1382.340 4.300 ;
        RECT 1383.500 2.890 1387.940 4.300 ;
        RECT 1389.100 2.890 1393.540 4.300 ;
        RECT 1394.700 2.890 1399.140 4.300 ;
        RECT 1400.300 2.890 1404.740 4.300 ;
        RECT 1405.900 2.890 1410.340 4.300 ;
        RECT 1411.500 2.890 1415.940 4.300 ;
        RECT 1417.100 2.890 1421.540 4.300 ;
        RECT 1422.700 2.890 1427.140 4.300 ;
        RECT 1428.300 2.890 1432.740 4.300 ;
        RECT 1433.900 2.890 1438.340 4.300 ;
        RECT 1439.500 2.890 1443.940 4.300 ;
        RECT 1445.100 2.890 1449.540 4.300 ;
        RECT 1450.700 2.890 1455.140 4.300 ;
        RECT 1456.300 2.890 1460.740 4.300 ;
        RECT 1461.900 2.890 1466.340 4.300 ;
        RECT 1467.500 2.890 1471.940 4.300 ;
        RECT 1473.100 2.890 1477.540 4.300 ;
        RECT 1478.700 2.890 1483.140 4.300 ;
        RECT 1484.300 2.890 1488.740 4.300 ;
        RECT 1489.900 2.890 1494.340 4.300 ;
        RECT 1495.500 2.890 1499.940 4.300 ;
        RECT 1501.100 2.890 1505.540 4.300 ;
        RECT 1506.700 2.890 1511.140 4.300 ;
        RECT 1512.300 2.890 1516.740 4.300 ;
        RECT 1517.900 2.890 1522.340 4.300 ;
        RECT 1523.500 2.890 1527.940 4.300 ;
        RECT 1529.100 2.890 1533.540 4.300 ;
        RECT 1534.700 2.890 1539.140 4.300 ;
        RECT 1540.300 2.890 1544.740 4.300 ;
        RECT 1545.900 2.890 1550.340 4.300 ;
        RECT 1551.500 2.890 1555.940 4.300 ;
        RECT 1557.100 2.890 1561.540 4.300 ;
        RECT 1562.700 2.890 1567.140 4.300 ;
        RECT 1568.300 2.890 1572.740 4.300 ;
        RECT 1573.900 2.890 1578.340 4.300 ;
        RECT 1579.500 2.890 1583.940 4.300 ;
        RECT 1585.100 2.890 1589.540 4.300 ;
        RECT 1590.700 2.890 1595.140 4.300 ;
        RECT 1596.300 2.890 1600.740 4.300 ;
        RECT 1601.900 2.890 1606.340 4.300 ;
        RECT 1607.500 2.890 1611.940 4.300 ;
        RECT 1613.100 2.890 1617.540 4.300 ;
        RECT 1618.700 2.890 1623.140 4.300 ;
        RECT 1624.300 2.890 1628.740 4.300 ;
        RECT 1629.900 2.890 1634.340 4.300 ;
        RECT 1635.500 2.890 1639.940 4.300 ;
        RECT 1641.100 2.890 1645.540 4.300 ;
        RECT 1646.700 2.890 1651.140 4.300 ;
        RECT 1652.300 2.890 1656.740 4.300 ;
        RECT 1657.900 2.890 1662.340 4.300 ;
        RECT 1663.500 2.890 1667.940 4.300 ;
        RECT 1669.100 2.890 1673.540 4.300 ;
        RECT 1674.700 2.890 1679.140 4.300 ;
        RECT 1680.300 2.890 1684.740 4.300 ;
        RECT 1685.900 2.890 1690.340 4.300 ;
        RECT 1691.500 2.890 1695.940 4.300 ;
        RECT 1697.100 2.890 1701.540 4.300 ;
        RECT 1702.700 2.890 1707.140 4.300 ;
        RECT 1708.300 2.890 1712.740 4.300 ;
        RECT 1713.900 2.890 1718.340 4.300 ;
        RECT 1719.500 2.890 1723.940 4.300 ;
        RECT 1725.100 2.890 1729.540 4.300 ;
        RECT 1730.700 2.890 1735.140 4.300 ;
        RECT 1736.300 2.890 1740.740 4.300 ;
        RECT 1741.900 2.890 1746.340 4.300 ;
        RECT 1747.500 2.890 1751.940 4.300 ;
        RECT 1753.100 2.890 1757.540 4.300 ;
        RECT 1758.700 2.890 1763.140 4.300 ;
        RECT 1764.300 2.890 1768.740 4.300 ;
        RECT 1769.900 2.890 1774.340 4.300 ;
        RECT 1775.500 2.890 1779.940 4.300 ;
        RECT 1781.100 2.890 1785.540 4.300 ;
        RECT 1786.700 2.890 1791.140 4.300 ;
        RECT 1792.300 2.890 1796.740 4.300 ;
        RECT 1797.900 2.890 1802.340 4.300 ;
        RECT 1803.500 2.890 1807.940 4.300 ;
        RECT 1809.100 2.890 1813.540 4.300 ;
        RECT 1814.700 2.890 1819.140 4.300 ;
        RECT 1820.300 2.890 1824.740 4.300 ;
        RECT 1825.900 2.890 1830.340 4.300 ;
        RECT 1831.500 2.890 1835.940 4.300 ;
        RECT 1837.100 2.890 1841.540 4.300 ;
        RECT 1842.700 2.890 1847.140 4.300 ;
        RECT 1848.300 2.890 1852.740 4.300 ;
        RECT 1853.900 2.890 1858.340 4.300 ;
        RECT 1859.500 2.890 1863.940 4.300 ;
        RECT 1865.100 2.890 1869.540 4.300 ;
        RECT 1870.700 2.890 1875.140 4.300 ;
        RECT 1876.300 2.890 1880.740 4.300 ;
        RECT 1881.900 2.890 1886.340 4.300 ;
        RECT 1887.500 2.890 1891.940 4.300 ;
        RECT 1893.100 2.890 1897.540 4.300 ;
        RECT 1898.700 2.890 1903.140 4.300 ;
        RECT 1904.300 2.890 1908.740 4.300 ;
        RECT 1909.900 2.890 1914.340 4.300 ;
        RECT 1915.500 2.890 1919.940 4.300 ;
        RECT 1921.100 2.890 1925.540 4.300 ;
        RECT 1926.700 2.890 1931.140 4.300 ;
        RECT 1932.300 2.890 1936.740 4.300 ;
        RECT 1937.900 2.890 1942.340 4.300 ;
        RECT 1943.500 2.890 1947.940 4.300 ;
        RECT 1949.100 2.890 1953.540 4.300 ;
        RECT 1954.700 2.890 1959.140 4.300 ;
        RECT 1960.300 2.890 1964.740 4.300 ;
        RECT 1965.900 2.890 1970.340 4.300 ;
        RECT 1971.500 2.890 1975.940 4.300 ;
        RECT 1977.100 2.890 1981.540 4.300 ;
        RECT 1982.700 2.890 1987.140 4.300 ;
        RECT 1988.300 2.890 1992.740 4.300 ;
        RECT 1993.900 2.890 1998.340 4.300 ;
        RECT 1999.500 2.890 2003.940 4.300 ;
        RECT 2005.100 2.890 2009.540 4.300 ;
        RECT 2010.700 2.890 2015.140 4.300 ;
        RECT 2016.300 2.890 2020.740 4.300 ;
        RECT 2021.900 2.890 2026.340 4.300 ;
        RECT 2027.500 2.890 2031.940 4.300 ;
        RECT 2033.100 2.890 2037.540 4.300 ;
        RECT 2038.700 2.890 2043.140 4.300 ;
        RECT 2044.300 2.890 2048.740 4.300 ;
        RECT 2049.900 2.890 2054.340 4.300 ;
        RECT 2055.500 2.890 2059.940 4.300 ;
        RECT 2061.100 2.890 2065.540 4.300 ;
        RECT 2066.700 2.890 2071.140 4.300 ;
        RECT 2072.300 2.890 2076.740 4.300 ;
        RECT 2077.900 2.890 2082.340 4.300 ;
        RECT 2083.500 2.890 2087.940 4.300 ;
        RECT 2089.100 2.890 2093.540 4.300 ;
        RECT 2094.700 2.890 2099.140 4.300 ;
        RECT 2100.300 2.890 2104.740 4.300 ;
        RECT 2105.900 2.890 2110.340 4.300 ;
        RECT 2111.500 2.890 2115.940 4.300 ;
        RECT 2117.100 2.890 2121.540 4.300 ;
        RECT 2122.700 2.890 2127.140 4.300 ;
        RECT 2128.300 2.890 2132.740 4.300 ;
        RECT 2133.900 2.890 2138.340 4.300 ;
        RECT 2139.500 2.890 2143.940 4.300 ;
        RECT 2145.100 2.890 2149.540 4.300 ;
        RECT 2150.700 2.890 2155.140 4.300 ;
        RECT 2156.300 2.890 2160.740 4.300 ;
        RECT 2161.900 2.890 2166.340 4.300 ;
        RECT 2167.500 2.890 2171.940 4.300 ;
        RECT 2173.100 2.890 2177.540 4.300 ;
        RECT 2178.700 2.890 2183.140 4.300 ;
        RECT 2184.300 2.890 2188.740 4.300 ;
        RECT 2189.900 2.890 2194.340 4.300 ;
        RECT 2195.500 2.890 2199.940 4.300 ;
        RECT 2201.100 2.890 2205.540 4.300 ;
        RECT 2206.700 2.890 2211.140 4.300 ;
        RECT 2212.300 2.890 2216.740 4.300 ;
        RECT 2217.900 2.890 2222.340 4.300 ;
        RECT 2223.500 2.890 2227.940 4.300 ;
        RECT 2229.100 2.890 2233.540 4.300 ;
        RECT 2234.700 2.890 2239.140 4.300 ;
        RECT 2240.300 2.890 2244.740 4.300 ;
        RECT 2245.900 2.890 2250.340 4.300 ;
        RECT 2251.500 2.890 2255.940 4.300 ;
        RECT 2257.100 2.890 2261.540 4.300 ;
        RECT 2262.700 2.890 2267.140 4.300 ;
        RECT 2268.300 2.890 2272.740 4.300 ;
        RECT 2273.900 2.890 2278.340 4.300 ;
        RECT 2279.500 2.890 2283.940 4.300 ;
        RECT 2285.100 2.890 2289.540 4.300 ;
        RECT 2290.700 2.890 2295.140 4.300 ;
        RECT 2296.300 2.890 2300.740 4.300 ;
        RECT 2301.900 2.890 2306.340 4.300 ;
        RECT 2307.500 2.890 2311.940 4.300 ;
        RECT 2313.100 2.890 2317.540 4.300 ;
        RECT 2318.700 2.890 2323.140 4.300 ;
        RECT 2324.300 2.890 2328.740 4.300 ;
        RECT 2329.900 2.890 2334.340 4.300 ;
        RECT 2335.500 2.890 2339.940 4.300 ;
        RECT 2341.100 2.890 2345.540 4.300 ;
        RECT 2346.700 2.890 2351.140 4.300 ;
        RECT 2352.300 2.890 2356.740 4.300 ;
        RECT 2357.900 2.890 2362.340 4.300 ;
        RECT 2363.500 2.890 2367.940 4.300 ;
        RECT 2369.100 2.890 2373.540 4.300 ;
        RECT 2374.700 2.890 2379.140 4.300 ;
        RECT 2380.300 2.890 2384.740 4.300 ;
        RECT 2385.900 2.890 2390.340 4.300 ;
        RECT 2391.500 2.890 2395.940 4.300 ;
        RECT 2397.100 2.890 2401.540 4.300 ;
        RECT 2402.700 2.890 2407.140 4.300 ;
        RECT 2408.300 2.890 2412.740 4.300 ;
        RECT 2413.900 2.890 2418.340 4.300 ;
        RECT 2419.500 2.890 2423.940 4.300 ;
        RECT 2425.100 2.890 2429.540 4.300 ;
        RECT 2430.700 2.890 2435.140 4.300 ;
        RECT 2436.300 2.890 2440.740 4.300 ;
        RECT 2441.900 2.890 2446.340 4.300 ;
        RECT 2447.500 2.890 2451.940 4.300 ;
        RECT 2453.100 2.890 2457.540 4.300 ;
        RECT 2458.700 2.890 2463.140 4.300 ;
        RECT 2464.300 2.890 2468.740 4.300 ;
        RECT 2469.900 2.890 2474.340 4.300 ;
        RECT 2475.500 2.890 2479.940 4.300 ;
        RECT 2481.100 2.890 2485.540 4.300 ;
        RECT 2486.700 2.890 2491.140 4.300 ;
        RECT 2492.300 2.890 2496.740 4.300 ;
        RECT 2497.900 2.890 2502.340 4.300 ;
        RECT 2503.500 2.890 2507.940 4.300 ;
        RECT 2509.100 2.890 2513.540 4.300 ;
        RECT 2514.700 2.890 2519.140 4.300 ;
        RECT 2520.300 2.890 2524.740 4.300 ;
        RECT 2525.900 2.890 2530.340 4.300 ;
        RECT 2531.500 2.890 2535.940 4.300 ;
        RECT 2537.100 2.890 2541.540 4.300 ;
        RECT 2542.700 2.890 2547.140 4.300 ;
        RECT 2548.300 2.890 2552.740 4.300 ;
        RECT 2553.900 2.890 2558.340 4.300 ;
        RECT 2559.500 2.890 2563.940 4.300 ;
        RECT 2565.100 2.890 2569.540 4.300 ;
        RECT 2570.700 2.890 2575.140 4.300 ;
        RECT 2576.300 2.890 2580.740 4.300 ;
        RECT 2581.900 2.890 2586.340 4.300 ;
        RECT 2587.500 2.890 2591.940 4.300 ;
        RECT 2593.100 2.890 2597.540 4.300 ;
        RECT 2598.700 2.890 2603.140 4.300 ;
        RECT 2604.300 2.890 2608.740 4.300 ;
        RECT 2609.900 2.890 2614.340 4.300 ;
        RECT 2615.500 2.890 2619.940 4.300 ;
        RECT 2621.100 2.890 2625.540 4.300 ;
        RECT 2626.700 2.890 2631.140 4.300 ;
        RECT 2632.300 2.890 2636.740 4.300 ;
        RECT 2637.900 2.890 2642.340 4.300 ;
        RECT 2643.500 2.890 2647.940 4.300 ;
        RECT 2649.100 2.890 2653.540 4.300 ;
        RECT 2654.700 2.890 2659.140 4.300 ;
        RECT 2660.300 2.890 2664.740 4.300 ;
        RECT 2665.900 2.890 2670.340 4.300 ;
        RECT 2671.500 2.890 2675.940 4.300 ;
        RECT 2677.100 2.890 2681.540 4.300 ;
        RECT 2682.700 2.890 2687.140 4.300 ;
        RECT 2688.300 2.890 2692.740 4.300 ;
        RECT 2693.900 2.890 2698.340 4.300 ;
        RECT 2699.500 2.890 2703.940 4.300 ;
        RECT 2705.100 2.890 2709.540 4.300 ;
        RECT 2710.700 2.890 2715.140 4.300 ;
        RECT 2716.300 2.890 2720.740 4.300 ;
        RECT 2721.900 2.890 2726.340 4.300 ;
        RECT 2727.500 2.890 2731.940 4.300 ;
        RECT 2733.100 2.890 2737.540 4.300 ;
        RECT 2738.700 2.890 2743.140 4.300 ;
        RECT 2744.300 2.890 2748.740 4.300 ;
        RECT 2749.900 2.890 2754.340 4.300 ;
        RECT 2755.500 2.890 2759.940 4.300 ;
        RECT 2761.100 2.890 2765.540 4.300 ;
        RECT 2766.700 2.890 2771.140 4.300 ;
        RECT 2772.300 2.890 2776.740 4.300 ;
        RECT 2777.900 2.890 2792.580 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 1717.820 2796.000 1740.620 ;
        RECT 4.300 1716.660 2795.700 1717.820 ;
        RECT 4.000 1645.020 2796.000 1716.660 ;
        RECT 4.300 1643.860 2795.700 1645.020 ;
        RECT 4.000 1572.220 2796.000 1643.860 ;
        RECT 4.300 1571.060 2795.700 1572.220 ;
        RECT 4.000 1499.420 2796.000 1571.060 ;
        RECT 4.300 1498.260 2795.700 1499.420 ;
        RECT 4.000 1426.620 2796.000 1498.260 ;
        RECT 4.300 1425.460 2795.700 1426.620 ;
        RECT 4.000 1353.820 2796.000 1425.460 ;
        RECT 4.300 1352.660 2795.700 1353.820 ;
        RECT 4.000 1281.020 2796.000 1352.660 ;
        RECT 4.300 1279.860 2795.700 1281.020 ;
        RECT 4.000 1208.220 2796.000 1279.860 ;
        RECT 4.300 1207.060 2795.700 1208.220 ;
        RECT 4.000 1135.420 2796.000 1207.060 ;
        RECT 4.300 1134.260 2795.700 1135.420 ;
        RECT 4.000 1062.620 2796.000 1134.260 ;
        RECT 4.300 1061.460 2795.700 1062.620 ;
        RECT 4.000 989.820 2796.000 1061.460 ;
        RECT 4.300 988.660 2795.700 989.820 ;
        RECT 4.000 917.020 2796.000 988.660 ;
        RECT 4.300 915.860 2795.700 917.020 ;
        RECT 4.000 844.220 2796.000 915.860 ;
        RECT 4.300 843.060 2795.700 844.220 ;
        RECT 4.000 771.420 2796.000 843.060 ;
        RECT 4.300 770.260 2795.700 771.420 ;
        RECT 4.000 698.620 2796.000 770.260 ;
        RECT 4.300 697.460 2795.700 698.620 ;
        RECT 4.000 625.820 2796.000 697.460 ;
        RECT 4.300 624.660 2795.700 625.820 ;
        RECT 4.000 553.020 2796.000 624.660 ;
        RECT 4.300 551.860 2795.700 553.020 ;
        RECT 4.000 480.220 2796.000 551.860 ;
        RECT 4.300 479.060 2795.700 480.220 ;
        RECT 4.000 407.420 2796.000 479.060 ;
        RECT 4.300 406.260 2795.700 407.420 ;
        RECT 4.000 334.620 2796.000 406.260 ;
        RECT 4.300 333.460 2795.700 334.620 ;
        RECT 4.000 261.820 2796.000 333.460 ;
        RECT 4.300 260.660 2795.700 261.820 ;
        RECT 4.000 189.020 2796.000 260.660 ;
        RECT 4.300 187.860 2795.700 189.020 ;
        RECT 4.000 116.220 2796.000 187.860 ;
        RECT 4.300 115.060 2795.700 116.220 ;
        RECT 4.000 43.420 2796.000 115.060 ;
        RECT 4.300 42.260 2795.700 43.420 ;
        RECT 4.000 2.940 2796.000 42.260 ;
      LAYER Metal4 ;
        RECT 775.740 15.080 789.940 41.350 ;
        RECT 792.140 15.080 866.740 41.350 ;
        RECT 868.940 15.080 943.540 41.350 ;
        RECT 945.740 15.080 1020.340 41.350 ;
        RECT 1022.540 15.080 1097.140 41.350 ;
        RECT 1099.340 15.080 1173.940 41.350 ;
        RECT 1176.140 15.080 1223.460 41.350 ;
        RECT 775.740 4.010 1223.460 15.080 ;
  END
END user_proj_example
END LIBRARY

