magic
tech gf180mcuC
magscale 1 5
timestamp 1688985070
<< obsm1 >>
rect 672 855 279328 174078
<< metal2 >>
rect 2184 0 2240 400
rect 2744 0 2800 400
rect 3304 0 3360 400
rect 3864 0 3920 400
rect 4424 0 4480 400
rect 4984 0 5040 400
rect 5544 0 5600 400
rect 6104 0 6160 400
rect 6664 0 6720 400
rect 7224 0 7280 400
rect 7784 0 7840 400
rect 8344 0 8400 400
rect 8904 0 8960 400
rect 9464 0 9520 400
rect 10024 0 10080 400
rect 10584 0 10640 400
rect 11144 0 11200 400
rect 11704 0 11760 400
rect 12264 0 12320 400
rect 12824 0 12880 400
rect 13384 0 13440 400
rect 13944 0 14000 400
rect 14504 0 14560 400
rect 15064 0 15120 400
rect 15624 0 15680 400
rect 16184 0 16240 400
rect 16744 0 16800 400
rect 17304 0 17360 400
rect 17864 0 17920 400
rect 18424 0 18480 400
rect 18984 0 19040 400
rect 19544 0 19600 400
rect 20104 0 20160 400
rect 20664 0 20720 400
rect 21224 0 21280 400
rect 21784 0 21840 400
rect 22344 0 22400 400
rect 22904 0 22960 400
rect 23464 0 23520 400
rect 24024 0 24080 400
rect 24584 0 24640 400
rect 25144 0 25200 400
rect 25704 0 25760 400
rect 26264 0 26320 400
rect 26824 0 26880 400
rect 27384 0 27440 400
rect 27944 0 28000 400
rect 28504 0 28560 400
rect 29064 0 29120 400
rect 29624 0 29680 400
rect 30184 0 30240 400
rect 30744 0 30800 400
rect 31304 0 31360 400
rect 31864 0 31920 400
rect 32424 0 32480 400
rect 32984 0 33040 400
rect 33544 0 33600 400
rect 34104 0 34160 400
rect 34664 0 34720 400
rect 35224 0 35280 400
rect 35784 0 35840 400
rect 36344 0 36400 400
rect 36904 0 36960 400
rect 37464 0 37520 400
rect 38024 0 38080 400
rect 38584 0 38640 400
rect 39144 0 39200 400
rect 39704 0 39760 400
rect 40264 0 40320 400
rect 40824 0 40880 400
rect 41384 0 41440 400
rect 41944 0 42000 400
rect 42504 0 42560 400
rect 43064 0 43120 400
rect 43624 0 43680 400
rect 44184 0 44240 400
rect 44744 0 44800 400
rect 45304 0 45360 400
rect 45864 0 45920 400
rect 46424 0 46480 400
rect 46984 0 47040 400
rect 47544 0 47600 400
rect 48104 0 48160 400
rect 48664 0 48720 400
rect 49224 0 49280 400
rect 49784 0 49840 400
rect 50344 0 50400 400
rect 50904 0 50960 400
rect 51464 0 51520 400
rect 52024 0 52080 400
rect 52584 0 52640 400
rect 53144 0 53200 400
rect 53704 0 53760 400
rect 54264 0 54320 400
rect 54824 0 54880 400
rect 55384 0 55440 400
rect 55944 0 56000 400
rect 56504 0 56560 400
rect 57064 0 57120 400
rect 57624 0 57680 400
rect 58184 0 58240 400
rect 58744 0 58800 400
rect 59304 0 59360 400
rect 59864 0 59920 400
rect 60424 0 60480 400
rect 60984 0 61040 400
rect 61544 0 61600 400
rect 62104 0 62160 400
rect 62664 0 62720 400
rect 63224 0 63280 400
rect 63784 0 63840 400
rect 64344 0 64400 400
rect 64904 0 64960 400
rect 65464 0 65520 400
rect 66024 0 66080 400
rect 66584 0 66640 400
rect 67144 0 67200 400
rect 67704 0 67760 400
rect 68264 0 68320 400
rect 68824 0 68880 400
rect 69384 0 69440 400
rect 69944 0 70000 400
rect 70504 0 70560 400
rect 71064 0 71120 400
rect 71624 0 71680 400
rect 72184 0 72240 400
rect 72744 0 72800 400
rect 73304 0 73360 400
rect 73864 0 73920 400
rect 74424 0 74480 400
rect 74984 0 75040 400
rect 75544 0 75600 400
rect 76104 0 76160 400
rect 76664 0 76720 400
rect 77224 0 77280 400
rect 77784 0 77840 400
rect 78344 0 78400 400
rect 78904 0 78960 400
rect 79464 0 79520 400
rect 80024 0 80080 400
rect 80584 0 80640 400
rect 81144 0 81200 400
rect 81704 0 81760 400
rect 82264 0 82320 400
rect 82824 0 82880 400
rect 83384 0 83440 400
rect 83944 0 84000 400
rect 84504 0 84560 400
rect 85064 0 85120 400
rect 85624 0 85680 400
rect 86184 0 86240 400
rect 86744 0 86800 400
rect 87304 0 87360 400
rect 87864 0 87920 400
rect 88424 0 88480 400
rect 88984 0 89040 400
rect 89544 0 89600 400
rect 90104 0 90160 400
rect 90664 0 90720 400
rect 91224 0 91280 400
rect 91784 0 91840 400
rect 92344 0 92400 400
rect 92904 0 92960 400
rect 93464 0 93520 400
rect 94024 0 94080 400
rect 94584 0 94640 400
rect 95144 0 95200 400
rect 95704 0 95760 400
rect 96264 0 96320 400
rect 96824 0 96880 400
rect 97384 0 97440 400
rect 97944 0 98000 400
rect 98504 0 98560 400
rect 99064 0 99120 400
rect 99624 0 99680 400
rect 100184 0 100240 400
rect 100744 0 100800 400
rect 101304 0 101360 400
rect 101864 0 101920 400
rect 102424 0 102480 400
rect 102984 0 103040 400
rect 103544 0 103600 400
rect 104104 0 104160 400
rect 104664 0 104720 400
rect 105224 0 105280 400
rect 105784 0 105840 400
rect 106344 0 106400 400
rect 106904 0 106960 400
rect 107464 0 107520 400
rect 108024 0 108080 400
rect 108584 0 108640 400
rect 109144 0 109200 400
rect 109704 0 109760 400
rect 110264 0 110320 400
rect 110824 0 110880 400
rect 111384 0 111440 400
rect 111944 0 112000 400
rect 112504 0 112560 400
rect 113064 0 113120 400
rect 113624 0 113680 400
rect 114184 0 114240 400
rect 114744 0 114800 400
rect 115304 0 115360 400
rect 115864 0 115920 400
rect 116424 0 116480 400
rect 116984 0 117040 400
rect 117544 0 117600 400
rect 118104 0 118160 400
rect 118664 0 118720 400
rect 119224 0 119280 400
rect 119784 0 119840 400
rect 120344 0 120400 400
rect 120904 0 120960 400
rect 121464 0 121520 400
rect 122024 0 122080 400
rect 122584 0 122640 400
rect 123144 0 123200 400
rect 123704 0 123760 400
rect 124264 0 124320 400
rect 124824 0 124880 400
rect 125384 0 125440 400
rect 125944 0 126000 400
rect 126504 0 126560 400
rect 127064 0 127120 400
rect 127624 0 127680 400
rect 128184 0 128240 400
rect 128744 0 128800 400
rect 129304 0 129360 400
rect 129864 0 129920 400
rect 130424 0 130480 400
rect 130984 0 131040 400
rect 131544 0 131600 400
rect 132104 0 132160 400
rect 132664 0 132720 400
rect 133224 0 133280 400
rect 133784 0 133840 400
rect 134344 0 134400 400
rect 134904 0 134960 400
rect 135464 0 135520 400
rect 136024 0 136080 400
rect 136584 0 136640 400
rect 137144 0 137200 400
rect 137704 0 137760 400
rect 138264 0 138320 400
rect 138824 0 138880 400
rect 139384 0 139440 400
rect 139944 0 140000 400
rect 140504 0 140560 400
rect 141064 0 141120 400
rect 141624 0 141680 400
rect 142184 0 142240 400
rect 142744 0 142800 400
rect 143304 0 143360 400
rect 143864 0 143920 400
rect 144424 0 144480 400
rect 144984 0 145040 400
rect 145544 0 145600 400
rect 146104 0 146160 400
rect 146664 0 146720 400
rect 147224 0 147280 400
rect 147784 0 147840 400
rect 148344 0 148400 400
rect 148904 0 148960 400
rect 149464 0 149520 400
rect 150024 0 150080 400
rect 150584 0 150640 400
rect 151144 0 151200 400
rect 151704 0 151760 400
rect 152264 0 152320 400
rect 152824 0 152880 400
rect 153384 0 153440 400
rect 153944 0 154000 400
rect 154504 0 154560 400
rect 155064 0 155120 400
rect 155624 0 155680 400
rect 156184 0 156240 400
rect 156744 0 156800 400
rect 157304 0 157360 400
rect 157864 0 157920 400
rect 158424 0 158480 400
rect 158984 0 159040 400
rect 159544 0 159600 400
rect 160104 0 160160 400
rect 160664 0 160720 400
rect 161224 0 161280 400
rect 161784 0 161840 400
rect 162344 0 162400 400
rect 162904 0 162960 400
rect 163464 0 163520 400
rect 164024 0 164080 400
rect 164584 0 164640 400
rect 165144 0 165200 400
rect 165704 0 165760 400
rect 166264 0 166320 400
rect 166824 0 166880 400
rect 167384 0 167440 400
rect 167944 0 168000 400
rect 168504 0 168560 400
rect 169064 0 169120 400
rect 169624 0 169680 400
rect 170184 0 170240 400
rect 170744 0 170800 400
rect 171304 0 171360 400
rect 171864 0 171920 400
rect 172424 0 172480 400
rect 172984 0 173040 400
rect 173544 0 173600 400
rect 174104 0 174160 400
rect 174664 0 174720 400
rect 175224 0 175280 400
rect 175784 0 175840 400
rect 176344 0 176400 400
rect 176904 0 176960 400
rect 177464 0 177520 400
rect 178024 0 178080 400
rect 178584 0 178640 400
rect 179144 0 179200 400
rect 179704 0 179760 400
rect 180264 0 180320 400
rect 180824 0 180880 400
rect 181384 0 181440 400
rect 181944 0 182000 400
rect 182504 0 182560 400
rect 183064 0 183120 400
rect 183624 0 183680 400
rect 184184 0 184240 400
rect 184744 0 184800 400
rect 185304 0 185360 400
rect 185864 0 185920 400
rect 186424 0 186480 400
rect 186984 0 187040 400
rect 187544 0 187600 400
rect 188104 0 188160 400
rect 188664 0 188720 400
rect 189224 0 189280 400
rect 189784 0 189840 400
rect 190344 0 190400 400
rect 190904 0 190960 400
rect 191464 0 191520 400
rect 192024 0 192080 400
rect 192584 0 192640 400
rect 193144 0 193200 400
rect 193704 0 193760 400
rect 194264 0 194320 400
rect 194824 0 194880 400
rect 195384 0 195440 400
rect 195944 0 196000 400
rect 196504 0 196560 400
rect 197064 0 197120 400
rect 197624 0 197680 400
rect 198184 0 198240 400
rect 198744 0 198800 400
rect 199304 0 199360 400
rect 199864 0 199920 400
rect 200424 0 200480 400
rect 200984 0 201040 400
rect 201544 0 201600 400
rect 202104 0 202160 400
rect 202664 0 202720 400
rect 203224 0 203280 400
rect 203784 0 203840 400
rect 204344 0 204400 400
rect 204904 0 204960 400
rect 205464 0 205520 400
rect 206024 0 206080 400
rect 206584 0 206640 400
rect 207144 0 207200 400
rect 207704 0 207760 400
rect 208264 0 208320 400
rect 208824 0 208880 400
rect 209384 0 209440 400
rect 209944 0 210000 400
rect 210504 0 210560 400
rect 211064 0 211120 400
rect 211624 0 211680 400
rect 212184 0 212240 400
rect 212744 0 212800 400
rect 213304 0 213360 400
rect 213864 0 213920 400
rect 214424 0 214480 400
rect 214984 0 215040 400
rect 215544 0 215600 400
rect 216104 0 216160 400
rect 216664 0 216720 400
rect 217224 0 217280 400
rect 217784 0 217840 400
rect 218344 0 218400 400
rect 218904 0 218960 400
rect 219464 0 219520 400
rect 220024 0 220080 400
rect 220584 0 220640 400
rect 221144 0 221200 400
rect 221704 0 221760 400
rect 222264 0 222320 400
rect 222824 0 222880 400
rect 223384 0 223440 400
rect 223944 0 224000 400
rect 224504 0 224560 400
rect 225064 0 225120 400
rect 225624 0 225680 400
rect 226184 0 226240 400
rect 226744 0 226800 400
rect 227304 0 227360 400
rect 227864 0 227920 400
rect 228424 0 228480 400
rect 228984 0 229040 400
rect 229544 0 229600 400
rect 230104 0 230160 400
rect 230664 0 230720 400
rect 231224 0 231280 400
rect 231784 0 231840 400
rect 232344 0 232400 400
rect 232904 0 232960 400
rect 233464 0 233520 400
rect 234024 0 234080 400
rect 234584 0 234640 400
rect 235144 0 235200 400
rect 235704 0 235760 400
rect 236264 0 236320 400
rect 236824 0 236880 400
rect 237384 0 237440 400
rect 237944 0 238000 400
rect 238504 0 238560 400
rect 239064 0 239120 400
rect 239624 0 239680 400
rect 240184 0 240240 400
rect 240744 0 240800 400
rect 241304 0 241360 400
rect 241864 0 241920 400
rect 242424 0 242480 400
rect 242984 0 243040 400
rect 243544 0 243600 400
rect 244104 0 244160 400
rect 244664 0 244720 400
rect 245224 0 245280 400
rect 245784 0 245840 400
rect 246344 0 246400 400
rect 246904 0 246960 400
rect 247464 0 247520 400
rect 248024 0 248080 400
rect 248584 0 248640 400
rect 249144 0 249200 400
rect 249704 0 249760 400
rect 250264 0 250320 400
rect 250824 0 250880 400
rect 251384 0 251440 400
rect 251944 0 252000 400
rect 252504 0 252560 400
rect 253064 0 253120 400
rect 253624 0 253680 400
rect 254184 0 254240 400
rect 254744 0 254800 400
rect 255304 0 255360 400
rect 255864 0 255920 400
rect 256424 0 256480 400
rect 256984 0 257040 400
rect 257544 0 257600 400
rect 258104 0 258160 400
rect 258664 0 258720 400
rect 259224 0 259280 400
rect 259784 0 259840 400
rect 260344 0 260400 400
rect 260904 0 260960 400
rect 261464 0 261520 400
rect 262024 0 262080 400
rect 262584 0 262640 400
rect 263144 0 263200 400
rect 263704 0 263760 400
rect 264264 0 264320 400
rect 264824 0 264880 400
rect 265384 0 265440 400
rect 265944 0 266000 400
rect 266504 0 266560 400
rect 267064 0 267120 400
rect 267624 0 267680 400
rect 268184 0 268240 400
rect 268744 0 268800 400
rect 269304 0 269360 400
rect 269864 0 269920 400
rect 270424 0 270480 400
rect 270984 0 271040 400
rect 271544 0 271600 400
rect 272104 0 272160 400
rect 272664 0 272720 400
rect 273224 0 273280 400
rect 273784 0 273840 400
rect 274344 0 274400 400
rect 274904 0 274960 400
rect 275464 0 275520 400
rect 276024 0 276080 400
rect 276584 0 276640 400
rect 277144 0 277200 400
rect 277704 0 277760 400
<< obsm2 >>
rect 462 430 279258 174067
rect 462 289 2154 430
rect 2270 289 2714 430
rect 2830 289 3274 430
rect 3390 289 3834 430
rect 3950 289 4394 430
rect 4510 289 4954 430
rect 5070 289 5514 430
rect 5630 289 6074 430
rect 6190 289 6634 430
rect 6750 289 7194 430
rect 7310 289 7754 430
rect 7870 289 8314 430
rect 8430 289 8874 430
rect 8990 289 9434 430
rect 9550 289 9994 430
rect 10110 289 10554 430
rect 10670 289 11114 430
rect 11230 289 11674 430
rect 11790 289 12234 430
rect 12350 289 12794 430
rect 12910 289 13354 430
rect 13470 289 13914 430
rect 14030 289 14474 430
rect 14590 289 15034 430
rect 15150 289 15594 430
rect 15710 289 16154 430
rect 16270 289 16714 430
rect 16830 289 17274 430
rect 17390 289 17834 430
rect 17950 289 18394 430
rect 18510 289 18954 430
rect 19070 289 19514 430
rect 19630 289 20074 430
rect 20190 289 20634 430
rect 20750 289 21194 430
rect 21310 289 21754 430
rect 21870 289 22314 430
rect 22430 289 22874 430
rect 22990 289 23434 430
rect 23550 289 23994 430
rect 24110 289 24554 430
rect 24670 289 25114 430
rect 25230 289 25674 430
rect 25790 289 26234 430
rect 26350 289 26794 430
rect 26910 289 27354 430
rect 27470 289 27914 430
rect 28030 289 28474 430
rect 28590 289 29034 430
rect 29150 289 29594 430
rect 29710 289 30154 430
rect 30270 289 30714 430
rect 30830 289 31274 430
rect 31390 289 31834 430
rect 31950 289 32394 430
rect 32510 289 32954 430
rect 33070 289 33514 430
rect 33630 289 34074 430
rect 34190 289 34634 430
rect 34750 289 35194 430
rect 35310 289 35754 430
rect 35870 289 36314 430
rect 36430 289 36874 430
rect 36990 289 37434 430
rect 37550 289 37994 430
rect 38110 289 38554 430
rect 38670 289 39114 430
rect 39230 289 39674 430
rect 39790 289 40234 430
rect 40350 289 40794 430
rect 40910 289 41354 430
rect 41470 289 41914 430
rect 42030 289 42474 430
rect 42590 289 43034 430
rect 43150 289 43594 430
rect 43710 289 44154 430
rect 44270 289 44714 430
rect 44830 289 45274 430
rect 45390 289 45834 430
rect 45950 289 46394 430
rect 46510 289 46954 430
rect 47070 289 47514 430
rect 47630 289 48074 430
rect 48190 289 48634 430
rect 48750 289 49194 430
rect 49310 289 49754 430
rect 49870 289 50314 430
rect 50430 289 50874 430
rect 50990 289 51434 430
rect 51550 289 51994 430
rect 52110 289 52554 430
rect 52670 289 53114 430
rect 53230 289 53674 430
rect 53790 289 54234 430
rect 54350 289 54794 430
rect 54910 289 55354 430
rect 55470 289 55914 430
rect 56030 289 56474 430
rect 56590 289 57034 430
rect 57150 289 57594 430
rect 57710 289 58154 430
rect 58270 289 58714 430
rect 58830 289 59274 430
rect 59390 289 59834 430
rect 59950 289 60394 430
rect 60510 289 60954 430
rect 61070 289 61514 430
rect 61630 289 62074 430
rect 62190 289 62634 430
rect 62750 289 63194 430
rect 63310 289 63754 430
rect 63870 289 64314 430
rect 64430 289 64874 430
rect 64990 289 65434 430
rect 65550 289 65994 430
rect 66110 289 66554 430
rect 66670 289 67114 430
rect 67230 289 67674 430
rect 67790 289 68234 430
rect 68350 289 68794 430
rect 68910 289 69354 430
rect 69470 289 69914 430
rect 70030 289 70474 430
rect 70590 289 71034 430
rect 71150 289 71594 430
rect 71710 289 72154 430
rect 72270 289 72714 430
rect 72830 289 73274 430
rect 73390 289 73834 430
rect 73950 289 74394 430
rect 74510 289 74954 430
rect 75070 289 75514 430
rect 75630 289 76074 430
rect 76190 289 76634 430
rect 76750 289 77194 430
rect 77310 289 77754 430
rect 77870 289 78314 430
rect 78430 289 78874 430
rect 78990 289 79434 430
rect 79550 289 79994 430
rect 80110 289 80554 430
rect 80670 289 81114 430
rect 81230 289 81674 430
rect 81790 289 82234 430
rect 82350 289 82794 430
rect 82910 289 83354 430
rect 83470 289 83914 430
rect 84030 289 84474 430
rect 84590 289 85034 430
rect 85150 289 85594 430
rect 85710 289 86154 430
rect 86270 289 86714 430
rect 86830 289 87274 430
rect 87390 289 87834 430
rect 87950 289 88394 430
rect 88510 289 88954 430
rect 89070 289 89514 430
rect 89630 289 90074 430
rect 90190 289 90634 430
rect 90750 289 91194 430
rect 91310 289 91754 430
rect 91870 289 92314 430
rect 92430 289 92874 430
rect 92990 289 93434 430
rect 93550 289 93994 430
rect 94110 289 94554 430
rect 94670 289 95114 430
rect 95230 289 95674 430
rect 95790 289 96234 430
rect 96350 289 96794 430
rect 96910 289 97354 430
rect 97470 289 97914 430
rect 98030 289 98474 430
rect 98590 289 99034 430
rect 99150 289 99594 430
rect 99710 289 100154 430
rect 100270 289 100714 430
rect 100830 289 101274 430
rect 101390 289 101834 430
rect 101950 289 102394 430
rect 102510 289 102954 430
rect 103070 289 103514 430
rect 103630 289 104074 430
rect 104190 289 104634 430
rect 104750 289 105194 430
rect 105310 289 105754 430
rect 105870 289 106314 430
rect 106430 289 106874 430
rect 106990 289 107434 430
rect 107550 289 107994 430
rect 108110 289 108554 430
rect 108670 289 109114 430
rect 109230 289 109674 430
rect 109790 289 110234 430
rect 110350 289 110794 430
rect 110910 289 111354 430
rect 111470 289 111914 430
rect 112030 289 112474 430
rect 112590 289 113034 430
rect 113150 289 113594 430
rect 113710 289 114154 430
rect 114270 289 114714 430
rect 114830 289 115274 430
rect 115390 289 115834 430
rect 115950 289 116394 430
rect 116510 289 116954 430
rect 117070 289 117514 430
rect 117630 289 118074 430
rect 118190 289 118634 430
rect 118750 289 119194 430
rect 119310 289 119754 430
rect 119870 289 120314 430
rect 120430 289 120874 430
rect 120990 289 121434 430
rect 121550 289 121994 430
rect 122110 289 122554 430
rect 122670 289 123114 430
rect 123230 289 123674 430
rect 123790 289 124234 430
rect 124350 289 124794 430
rect 124910 289 125354 430
rect 125470 289 125914 430
rect 126030 289 126474 430
rect 126590 289 127034 430
rect 127150 289 127594 430
rect 127710 289 128154 430
rect 128270 289 128714 430
rect 128830 289 129274 430
rect 129390 289 129834 430
rect 129950 289 130394 430
rect 130510 289 130954 430
rect 131070 289 131514 430
rect 131630 289 132074 430
rect 132190 289 132634 430
rect 132750 289 133194 430
rect 133310 289 133754 430
rect 133870 289 134314 430
rect 134430 289 134874 430
rect 134990 289 135434 430
rect 135550 289 135994 430
rect 136110 289 136554 430
rect 136670 289 137114 430
rect 137230 289 137674 430
rect 137790 289 138234 430
rect 138350 289 138794 430
rect 138910 289 139354 430
rect 139470 289 139914 430
rect 140030 289 140474 430
rect 140590 289 141034 430
rect 141150 289 141594 430
rect 141710 289 142154 430
rect 142270 289 142714 430
rect 142830 289 143274 430
rect 143390 289 143834 430
rect 143950 289 144394 430
rect 144510 289 144954 430
rect 145070 289 145514 430
rect 145630 289 146074 430
rect 146190 289 146634 430
rect 146750 289 147194 430
rect 147310 289 147754 430
rect 147870 289 148314 430
rect 148430 289 148874 430
rect 148990 289 149434 430
rect 149550 289 149994 430
rect 150110 289 150554 430
rect 150670 289 151114 430
rect 151230 289 151674 430
rect 151790 289 152234 430
rect 152350 289 152794 430
rect 152910 289 153354 430
rect 153470 289 153914 430
rect 154030 289 154474 430
rect 154590 289 155034 430
rect 155150 289 155594 430
rect 155710 289 156154 430
rect 156270 289 156714 430
rect 156830 289 157274 430
rect 157390 289 157834 430
rect 157950 289 158394 430
rect 158510 289 158954 430
rect 159070 289 159514 430
rect 159630 289 160074 430
rect 160190 289 160634 430
rect 160750 289 161194 430
rect 161310 289 161754 430
rect 161870 289 162314 430
rect 162430 289 162874 430
rect 162990 289 163434 430
rect 163550 289 163994 430
rect 164110 289 164554 430
rect 164670 289 165114 430
rect 165230 289 165674 430
rect 165790 289 166234 430
rect 166350 289 166794 430
rect 166910 289 167354 430
rect 167470 289 167914 430
rect 168030 289 168474 430
rect 168590 289 169034 430
rect 169150 289 169594 430
rect 169710 289 170154 430
rect 170270 289 170714 430
rect 170830 289 171274 430
rect 171390 289 171834 430
rect 171950 289 172394 430
rect 172510 289 172954 430
rect 173070 289 173514 430
rect 173630 289 174074 430
rect 174190 289 174634 430
rect 174750 289 175194 430
rect 175310 289 175754 430
rect 175870 289 176314 430
rect 176430 289 176874 430
rect 176990 289 177434 430
rect 177550 289 177994 430
rect 178110 289 178554 430
rect 178670 289 179114 430
rect 179230 289 179674 430
rect 179790 289 180234 430
rect 180350 289 180794 430
rect 180910 289 181354 430
rect 181470 289 181914 430
rect 182030 289 182474 430
rect 182590 289 183034 430
rect 183150 289 183594 430
rect 183710 289 184154 430
rect 184270 289 184714 430
rect 184830 289 185274 430
rect 185390 289 185834 430
rect 185950 289 186394 430
rect 186510 289 186954 430
rect 187070 289 187514 430
rect 187630 289 188074 430
rect 188190 289 188634 430
rect 188750 289 189194 430
rect 189310 289 189754 430
rect 189870 289 190314 430
rect 190430 289 190874 430
rect 190990 289 191434 430
rect 191550 289 191994 430
rect 192110 289 192554 430
rect 192670 289 193114 430
rect 193230 289 193674 430
rect 193790 289 194234 430
rect 194350 289 194794 430
rect 194910 289 195354 430
rect 195470 289 195914 430
rect 196030 289 196474 430
rect 196590 289 197034 430
rect 197150 289 197594 430
rect 197710 289 198154 430
rect 198270 289 198714 430
rect 198830 289 199274 430
rect 199390 289 199834 430
rect 199950 289 200394 430
rect 200510 289 200954 430
rect 201070 289 201514 430
rect 201630 289 202074 430
rect 202190 289 202634 430
rect 202750 289 203194 430
rect 203310 289 203754 430
rect 203870 289 204314 430
rect 204430 289 204874 430
rect 204990 289 205434 430
rect 205550 289 205994 430
rect 206110 289 206554 430
rect 206670 289 207114 430
rect 207230 289 207674 430
rect 207790 289 208234 430
rect 208350 289 208794 430
rect 208910 289 209354 430
rect 209470 289 209914 430
rect 210030 289 210474 430
rect 210590 289 211034 430
rect 211150 289 211594 430
rect 211710 289 212154 430
rect 212270 289 212714 430
rect 212830 289 213274 430
rect 213390 289 213834 430
rect 213950 289 214394 430
rect 214510 289 214954 430
rect 215070 289 215514 430
rect 215630 289 216074 430
rect 216190 289 216634 430
rect 216750 289 217194 430
rect 217310 289 217754 430
rect 217870 289 218314 430
rect 218430 289 218874 430
rect 218990 289 219434 430
rect 219550 289 219994 430
rect 220110 289 220554 430
rect 220670 289 221114 430
rect 221230 289 221674 430
rect 221790 289 222234 430
rect 222350 289 222794 430
rect 222910 289 223354 430
rect 223470 289 223914 430
rect 224030 289 224474 430
rect 224590 289 225034 430
rect 225150 289 225594 430
rect 225710 289 226154 430
rect 226270 289 226714 430
rect 226830 289 227274 430
rect 227390 289 227834 430
rect 227950 289 228394 430
rect 228510 289 228954 430
rect 229070 289 229514 430
rect 229630 289 230074 430
rect 230190 289 230634 430
rect 230750 289 231194 430
rect 231310 289 231754 430
rect 231870 289 232314 430
rect 232430 289 232874 430
rect 232990 289 233434 430
rect 233550 289 233994 430
rect 234110 289 234554 430
rect 234670 289 235114 430
rect 235230 289 235674 430
rect 235790 289 236234 430
rect 236350 289 236794 430
rect 236910 289 237354 430
rect 237470 289 237914 430
rect 238030 289 238474 430
rect 238590 289 239034 430
rect 239150 289 239594 430
rect 239710 289 240154 430
rect 240270 289 240714 430
rect 240830 289 241274 430
rect 241390 289 241834 430
rect 241950 289 242394 430
rect 242510 289 242954 430
rect 243070 289 243514 430
rect 243630 289 244074 430
rect 244190 289 244634 430
rect 244750 289 245194 430
rect 245310 289 245754 430
rect 245870 289 246314 430
rect 246430 289 246874 430
rect 246990 289 247434 430
rect 247550 289 247994 430
rect 248110 289 248554 430
rect 248670 289 249114 430
rect 249230 289 249674 430
rect 249790 289 250234 430
rect 250350 289 250794 430
rect 250910 289 251354 430
rect 251470 289 251914 430
rect 252030 289 252474 430
rect 252590 289 253034 430
rect 253150 289 253594 430
rect 253710 289 254154 430
rect 254270 289 254714 430
rect 254830 289 255274 430
rect 255390 289 255834 430
rect 255950 289 256394 430
rect 256510 289 256954 430
rect 257070 289 257514 430
rect 257630 289 258074 430
rect 258190 289 258634 430
rect 258750 289 259194 430
rect 259310 289 259754 430
rect 259870 289 260314 430
rect 260430 289 260874 430
rect 260990 289 261434 430
rect 261550 289 261994 430
rect 262110 289 262554 430
rect 262670 289 263114 430
rect 263230 289 263674 430
rect 263790 289 264234 430
rect 264350 289 264794 430
rect 264910 289 265354 430
rect 265470 289 265914 430
rect 266030 289 266474 430
rect 266590 289 267034 430
rect 267150 289 267594 430
rect 267710 289 268154 430
rect 268270 289 268714 430
rect 268830 289 269274 430
rect 269390 289 269834 430
rect 269950 289 270394 430
rect 270510 289 270954 430
rect 271070 289 271514 430
rect 271630 289 272074 430
rect 272190 289 272634 430
rect 272750 289 273194 430
rect 273310 289 273754 430
rect 273870 289 274314 430
rect 274430 289 274874 430
rect 274990 289 275434 430
rect 275550 289 275994 430
rect 276110 289 276554 430
rect 276670 289 277114 430
rect 277230 289 277674 430
rect 277790 289 279258 430
<< metal3 >>
rect 0 171696 400 171752
rect 279600 171696 280000 171752
rect 0 164416 400 164472
rect 279600 164416 280000 164472
rect 0 157136 400 157192
rect 279600 157136 280000 157192
rect 0 149856 400 149912
rect 279600 149856 280000 149912
rect 0 142576 400 142632
rect 279600 142576 280000 142632
rect 0 135296 400 135352
rect 279600 135296 280000 135352
rect 0 128016 400 128072
rect 279600 128016 280000 128072
rect 0 120736 400 120792
rect 279600 120736 280000 120792
rect 0 113456 400 113512
rect 279600 113456 280000 113512
rect 0 106176 400 106232
rect 279600 106176 280000 106232
rect 0 98896 400 98952
rect 279600 98896 280000 98952
rect 0 91616 400 91672
rect 279600 91616 280000 91672
rect 0 84336 400 84392
rect 279600 84336 280000 84392
rect 0 77056 400 77112
rect 279600 77056 280000 77112
rect 0 69776 400 69832
rect 279600 69776 280000 69832
rect 0 62496 400 62552
rect 279600 62496 280000 62552
rect 0 55216 400 55272
rect 279600 55216 280000 55272
rect 0 47936 400 47992
rect 279600 47936 280000 47992
rect 0 40656 400 40712
rect 279600 40656 280000 40712
rect 0 33376 400 33432
rect 279600 33376 280000 33432
rect 0 26096 400 26152
rect 279600 26096 280000 26152
rect 0 18816 400 18872
rect 279600 18816 280000 18872
rect 0 11536 400 11592
rect 279600 11536 280000 11592
rect 0 4256 400 4312
rect 279600 4256 280000 4312
<< obsm3 >>
rect 400 171782 279600 174062
rect 430 171666 279570 171782
rect 400 164502 279600 171666
rect 430 164386 279570 164502
rect 400 157222 279600 164386
rect 430 157106 279570 157222
rect 400 149942 279600 157106
rect 430 149826 279570 149942
rect 400 142662 279600 149826
rect 430 142546 279570 142662
rect 400 135382 279600 142546
rect 430 135266 279570 135382
rect 400 128102 279600 135266
rect 430 127986 279570 128102
rect 400 120822 279600 127986
rect 430 120706 279570 120822
rect 400 113542 279600 120706
rect 430 113426 279570 113542
rect 400 106262 279600 113426
rect 430 106146 279570 106262
rect 400 98982 279600 106146
rect 430 98866 279570 98982
rect 400 91702 279600 98866
rect 430 91586 279570 91702
rect 400 84422 279600 91586
rect 430 84306 279570 84422
rect 400 77142 279600 84306
rect 430 77026 279570 77142
rect 400 69862 279600 77026
rect 430 69746 279570 69862
rect 400 62582 279600 69746
rect 430 62466 279570 62582
rect 400 55302 279600 62466
rect 430 55186 279570 55302
rect 400 48022 279600 55186
rect 430 47906 279570 48022
rect 400 40742 279600 47906
rect 430 40626 279570 40742
rect 400 33462 279600 40626
rect 430 33346 279570 33462
rect 400 26182 279600 33346
rect 430 26066 279570 26182
rect 400 18902 279600 26066
rect 430 18786 279570 18902
rect 400 11622 279600 18786
rect 430 11506 279570 11622
rect 400 4342 279600 11506
rect 430 4226 279570 4342
rect 400 294 279600 4226
<< metal4 >>
rect 2224 1538 2384 174078
rect 9904 1538 10064 174078
rect 17584 1538 17744 174078
rect 25264 1538 25424 174078
rect 32944 1538 33104 174078
rect 40624 1538 40784 174078
rect 48304 1538 48464 174078
rect 55984 1538 56144 174078
rect 63664 1538 63824 174078
rect 71344 1538 71504 174078
rect 79024 1538 79184 174078
rect 86704 1538 86864 174078
rect 94384 1538 94544 174078
rect 102064 1538 102224 174078
rect 109744 1538 109904 174078
rect 117424 1538 117584 174078
rect 125104 1538 125264 174078
rect 132784 1538 132944 174078
rect 140464 1538 140624 174078
rect 148144 1538 148304 174078
rect 155824 1538 155984 174078
rect 163504 1538 163664 174078
rect 171184 1538 171344 174078
rect 178864 1538 179024 174078
rect 186544 1538 186704 174078
rect 194224 1538 194384 174078
rect 201904 1538 202064 174078
rect 209584 1538 209744 174078
rect 217264 1538 217424 174078
rect 224944 1538 225104 174078
rect 232624 1538 232784 174078
rect 240304 1538 240464 174078
rect 247984 1538 248144 174078
rect 255664 1538 255824 174078
rect 263344 1538 263504 174078
rect 271024 1538 271184 174078
rect 278704 1538 278864 174078
<< obsm4 >>
rect 77574 1508 78994 4135
rect 79214 1508 86674 4135
rect 86894 1508 94354 4135
rect 94574 1508 102034 4135
rect 102254 1508 109714 4135
rect 109934 1508 117394 4135
rect 117614 1508 122346 4135
rect 77574 401 122346 1508
<< labels >>
rlabel metal3 s 279600 4256 280000 4312 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 128016 400 128072 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 106176 400 106232 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 84336 400 84392 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 0 62496 400 62552 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 0 40656 400 40712 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 18816 400 18872 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 279600 26096 280000 26152 6 io_in[1]
port 8 nsew signal input
rlabel metal3 s 279600 47936 280000 47992 6 io_in[2]
port 9 nsew signal input
rlabel metal3 s 279600 69776 280000 69832 6 io_in[3]
port 10 nsew signal input
rlabel metal3 s 279600 91616 280000 91672 6 io_in[4]
port 11 nsew signal input
rlabel metal3 s 279600 113456 280000 113512 6 io_in[5]
port 12 nsew signal input
rlabel metal3 s 279600 135296 280000 135352 6 io_in[6]
port 13 nsew signal input
rlabel metal3 s 279600 157136 280000 157192 6 io_in[7]
port 14 nsew signal input
rlabel metal3 s 0 171696 400 171752 6 io_in[8]
port 15 nsew signal input
rlabel metal3 s 0 149856 400 149912 6 io_in[9]
port 16 nsew signal input
rlabel metal3 s 279600 18816 280000 18872 6 io_oeb[0]
port 17 nsew signal output
rlabel metal3 s 0 113456 400 113512 6 io_oeb[10]
port 18 nsew signal output
rlabel metal3 s 0 91616 400 91672 6 io_oeb[11]
port 19 nsew signal output
rlabel metal3 s 0 69776 400 69832 6 io_oeb[12]
port 20 nsew signal output
rlabel metal3 s 0 47936 400 47992 6 io_oeb[13]
port 21 nsew signal output
rlabel metal3 s 0 26096 400 26152 6 io_oeb[14]
port 22 nsew signal output
rlabel metal3 s 0 4256 400 4312 6 io_oeb[15]
port 23 nsew signal output
rlabel metal3 s 279600 40656 280000 40712 6 io_oeb[1]
port 24 nsew signal output
rlabel metal3 s 279600 62496 280000 62552 6 io_oeb[2]
port 25 nsew signal output
rlabel metal3 s 279600 84336 280000 84392 6 io_oeb[3]
port 26 nsew signal output
rlabel metal3 s 279600 106176 280000 106232 6 io_oeb[4]
port 27 nsew signal output
rlabel metal3 s 279600 128016 280000 128072 6 io_oeb[5]
port 28 nsew signal output
rlabel metal3 s 279600 149856 280000 149912 6 io_oeb[6]
port 29 nsew signal output
rlabel metal3 s 279600 171696 280000 171752 6 io_oeb[7]
port 30 nsew signal output
rlabel metal3 s 0 157136 400 157192 6 io_oeb[8]
port 31 nsew signal output
rlabel metal3 s 0 135296 400 135352 6 io_oeb[9]
port 32 nsew signal output
rlabel metal3 s 279600 11536 280000 11592 6 io_out[0]
port 33 nsew signal output
rlabel metal3 s 0 120736 400 120792 6 io_out[10]
port 34 nsew signal output
rlabel metal3 s 0 98896 400 98952 6 io_out[11]
port 35 nsew signal output
rlabel metal3 s 0 77056 400 77112 6 io_out[12]
port 36 nsew signal output
rlabel metal3 s 0 55216 400 55272 6 io_out[13]
port 37 nsew signal output
rlabel metal3 s 0 33376 400 33432 6 io_out[14]
port 38 nsew signal output
rlabel metal3 s 0 11536 400 11592 6 io_out[15]
port 39 nsew signal output
rlabel metal3 s 279600 33376 280000 33432 6 io_out[1]
port 40 nsew signal output
rlabel metal3 s 279600 55216 280000 55272 6 io_out[2]
port 41 nsew signal output
rlabel metal3 s 279600 77056 280000 77112 6 io_out[3]
port 42 nsew signal output
rlabel metal3 s 279600 98896 280000 98952 6 io_out[4]
port 43 nsew signal output
rlabel metal3 s 279600 120736 280000 120792 6 io_out[5]
port 44 nsew signal output
rlabel metal3 s 279600 142576 280000 142632 6 io_out[6]
port 45 nsew signal output
rlabel metal3 s 279600 164416 280000 164472 6 io_out[7]
port 46 nsew signal output
rlabel metal3 s 0 164416 400 164472 6 io_out[8]
port 47 nsew signal output
rlabel metal3 s 0 142576 400 142632 6 io_out[9]
port 48 nsew signal output
rlabel metal2 s 276584 0 276640 400 6 irq[0]
port 49 nsew signal output
rlabel metal2 s 277144 0 277200 400 6 irq[1]
port 50 nsew signal output
rlabel metal2 s 277704 0 277760 400 6 irq[2]
port 51 nsew signal output
rlabel metal2 s 61544 0 61600 400 6 la_data_in[0]
port 52 nsew signal input
rlabel metal2 s 229544 0 229600 400 6 la_data_in[100]
port 53 nsew signal input
rlabel metal2 s 231224 0 231280 400 6 la_data_in[101]
port 54 nsew signal input
rlabel metal2 s 232904 0 232960 400 6 la_data_in[102]
port 55 nsew signal input
rlabel metal2 s 234584 0 234640 400 6 la_data_in[103]
port 56 nsew signal input
rlabel metal2 s 236264 0 236320 400 6 la_data_in[104]
port 57 nsew signal input
rlabel metal2 s 237944 0 238000 400 6 la_data_in[105]
port 58 nsew signal input
rlabel metal2 s 239624 0 239680 400 6 la_data_in[106]
port 59 nsew signal input
rlabel metal2 s 241304 0 241360 400 6 la_data_in[107]
port 60 nsew signal input
rlabel metal2 s 242984 0 243040 400 6 la_data_in[108]
port 61 nsew signal input
rlabel metal2 s 244664 0 244720 400 6 la_data_in[109]
port 62 nsew signal input
rlabel metal2 s 78344 0 78400 400 6 la_data_in[10]
port 63 nsew signal input
rlabel metal2 s 246344 0 246400 400 6 la_data_in[110]
port 64 nsew signal input
rlabel metal2 s 248024 0 248080 400 6 la_data_in[111]
port 65 nsew signal input
rlabel metal2 s 249704 0 249760 400 6 la_data_in[112]
port 66 nsew signal input
rlabel metal2 s 251384 0 251440 400 6 la_data_in[113]
port 67 nsew signal input
rlabel metal2 s 253064 0 253120 400 6 la_data_in[114]
port 68 nsew signal input
rlabel metal2 s 254744 0 254800 400 6 la_data_in[115]
port 69 nsew signal input
rlabel metal2 s 256424 0 256480 400 6 la_data_in[116]
port 70 nsew signal input
rlabel metal2 s 258104 0 258160 400 6 la_data_in[117]
port 71 nsew signal input
rlabel metal2 s 259784 0 259840 400 6 la_data_in[118]
port 72 nsew signal input
rlabel metal2 s 261464 0 261520 400 6 la_data_in[119]
port 73 nsew signal input
rlabel metal2 s 80024 0 80080 400 6 la_data_in[11]
port 74 nsew signal input
rlabel metal2 s 263144 0 263200 400 6 la_data_in[120]
port 75 nsew signal input
rlabel metal2 s 264824 0 264880 400 6 la_data_in[121]
port 76 nsew signal input
rlabel metal2 s 266504 0 266560 400 6 la_data_in[122]
port 77 nsew signal input
rlabel metal2 s 268184 0 268240 400 6 la_data_in[123]
port 78 nsew signal input
rlabel metal2 s 269864 0 269920 400 6 la_data_in[124]
port 79 nsew signal input
rlabel metal2 s 271544 0 271600 400 6 la_data_in[125]
port 80 nsew signal input
rlabel metal2 s 273224 0 273280 400 6 la_data_in[126]
port 81 nsew signal input
rlabel metal2 s 274904 0 274960 400 6 la_data_in[127]
port 82 nsew signal input
rlabel metal2 s 81704 0 81760 400 6 la_data_in[12]
port 83 nsew signal input
rlabel metal2 s 83384 0 83440 400 6 la_data_in[13]
port 84 nsew signal input
rlabel metal2 s 85064 0 85120 400 6 la_data_in[14]
port 85 nsew signal input
rlabel metal2 s 86744 0 86800 400 6 la_data_in[15]
port 86 nsew signal input
rlabel metal2 s 88424 0 88480 400 6 la_data_in[16]
port 87 nsew signal input
rlabel metal2 s 90104 0 90160 400 6 la_data_in[17]
port 88 nsew signal input
rlabel metal2 s 91784 0 91840 400 6 la_data_in[18]
port 89 nsew signal input
rlabel metal2 s 93464 0 93520 400 6 la_data_in[19]
port 90 nsew signal input
rlabel metal2 s 63224 0 63280 400 6 la_data_in[1]
port 91 nsew signal input
rlabel metal2 s 95144 0 95200 400 6 la_data_in[20]
port 92 nsew signal input
rlabel metal2 s 96824 0 96880 400 6 la_data_in[21]
port 93 nsew signal input
rlabel metal2 s 98504 0 98560 400 6 la_data_in[22]
port 94 nsew signal input
rlabel metal2 s 100184 0 100240 400 6 la_data_in[23]
port 95 nsew signal input
rlabel metal2 s 101864 0 101920 400 6 la_data_in[24]
port 96 nsew signal input
rlabel metal2 s 103544 0 103600 400 6 la_data_in[25]
port 97 nsew signal input
rlabel metal2 s 105224 0 105280 400 6 la_data_in[26]
port 98 nsew signal input
rlabel metal2 s 106904 0 106960 400 6 la_data_in[27]
port 99 nsew signal input
rlabel metal2 s 108584 0 108640 400 6 la_data_in[28]
port 100 nsew signal input
rlabel metal2 s 110264 0 110320 400 6 la_data_in[29]
port 101 nsew signal input
rlabel metal2 s 64904 0 64960 400 6 la_data_in[2]
port 102 nsew signal input
rlabel metal2 s 111944 0 112000 400 6 la_data_in[30]
port 103 nsew signal input
rlabel metal2 s 113624 0 113680 400 6 la_data_in[31]
port 104 nsew signal input
rlabel metal2 s 115304 0 115360 400 6 la_data_in[32]
port 105 nsew signal input
rlabel metal2 s 116984 0 117040 400 6 la_data_in[33]
port 106 nsew signal input
rlabel metal2 s 118664 0 118720 400 6 la_data_in[34]
port 107 nsew signal input
rlabel metal2 s 120344 0 120400 400 6 la_data_in[35]
port 108 nsew signal input
rlabel metal2 s 122024 0 122080 400 6 la_data_in[36]
port 109 nsew signal input
rlabel metal2 s 123704 0 123760 400 6 la_data_in[37]
port 110 nsew signal input
rlabel metal2 s 125384 0 125440 400 6 la_data_in[38]
port 111 nsew signal input
rlabel metal2 s 127064 0 127120 400 6 la_data_in[39]
port 112 nsew signal input
rlabel metal2 s 66584 0 66640 400 6 la_data_in[3]
port 113 nsew signal input
rlabel metal2 s 128744 0 128800 400 6 la_data_in[40]
port 114 nsew signal input
rlabel metal2 s 130424 0 130480 400 6 la_data_in[41]
port 115 nsew signal input
rlabel metal2 s 132104 0 132160 400 6 la_data_in[42]
port 116 nsew signal input
rlabel metal2 s 133784 0 133840 400 6 la_data_in[43]
port 117 nsew signal input
rlabel metal2 s 135464 0 135520 400 6 la_data_in[44]
port 118 nsew signal input
rlabel metal2 s 137144 0 137200 400 6 la_data_in[45]
port 119 nsew signal input
rlabel metal2 s 138824 0 138880 400 6 la_data_in[46]
port 120 nsew signal input
rlabel metal2 s 140504 0 140560 400 6 la_data_in[47]
port 121 nsew signal input
rlabel metal2 s 142184 0 142240 400 6 la_data_in[48]
port 122 nsew signal input
rlabel metal2 s 143864 0 143920 400 6 la_data_in[49]
port 123 nsew signal input
rlabel metal2 s 68264 0 68320 400 6 la_data_in[4]
port 124 nsew signal input
rlabel metal2 s 145544 0 145600 400 6 la_data_in[50]
port 125 nsew signal input
rlabel metal2 s 147224 0 147280 400 6 la_data_in[51]
port 126 nsew signal input
rlabel metal2 s 148904 0 148960 400 6 la_data_in[52]
port 127 nsew signal input
rlabel metal2 s 150584 0 150640 400 6 la_data_in[53]
port 128 nsew signal input
rlabel metal2 s 152264 0 152320 400 6 la_data_in[54]
port 129 nsew signal input
rlabel metal2 s 153944 0 154000 400 6 la_data_in[55]
port 130 nsew signal input
rlabel metal2 s 155624 0 155680 400 6 la_data_in[56]
port 131 nsew signal input
rlabel metal2 s 157304 0 157360 400 6 la_data_in[57]
port 132 nsew signal input
rlabel metal2 s 158984 0 159040 400 6 la_data_in[58]
port 133 nsew signal input
rlabel metal2 s 160664 0 160720 400 6 la_data_in[59]
port 134 nsew signal input
rlabel metal2 s 69944 0 70000 400 6 la_data_in[5]
port 135 nsew signal input
rlabel metal2 s 162344 0 162400 400 6 la_data_in[60]
port 136 nsew signal input
rlabel metal2 s 164024 0 164080 400 6 la_data_in[61]
port 137 nsew signal input
rlabel metal2 s 165704 0 165760 400 6 la_data_in[62]
port 138 nsew signal input
rlabel metal2 s 167384 0 167440 400 6 la_data_in[63]
port 139 nsew signal input
rlabel metal2 s 169064 0 169120 400 6 la_data_in[64]
port 140 nsew signal input
rlabel metal2 s 170744 0 170800 400 6 la_data_in[65]
port 141 nsew signal input
rlabel metal2 s 172424 0 172480 400 6 la_data_in[66]
port 142 nsew signal input
rlabel metal2 s 174104 0 174160 400 6 la_data_in[67]
port 143 nsew signal input
rlabel metal2 s 175784 0 175840 400 6 la_data_in[68]
port 144 nsew signal input
rlabel metal2 s 177464 0 177520 400 6 la_data_in[69]
port 145 nsew signal input
rlabel metal2 s 71624 0 71680 400 6 la_data_in[6]
port 146 nsew signal input
rlabel metal2 s 179144 0 179200 400 6 la_data_in[70]
port 147 nsew signal input
rlabel metal2 s 180824 0 180880 400 6 la_data_in[71]
port 148 nsew signal input
rlabel metal2 s 182504 0 182560 400 6 la_data_in[72]
port 149 nsew signal input
rlabel metal2 s 184184 0 184240 400 6 la_data_in[73]
port 150 nsew signal input
rlabel metal2 s 185864 0 185920 400 6 la_data_in[74]
port 151 nsew signal input
rlabel metal2 s 187544 0 187600 400 6 la_data_in[75]
port 152 nsew signal input
rlabel metal2 s 189224 0 189280 400 6 la_data_in[76]
port 153 nsew signal input
rlabel metal2 s 190904 0 190960 400 6 la_data_in[77]
port 154 nsew signal input
rlabel metal2 s 192584 0 192640 400 6 la_data_in[78]
port 155 nsew signal input
rlabel metal2 s 194264 0 194320 400 6 la_data_in[79]
port 156 nsew signal input
rlabel metal2 s 73304 0 73360 400 6 la_data_in[7]
port 157 nsew signal input
rlabel metal2 s 195944 0 196000 400 6 la_data_in[80]
port 158 nsew signal input
rlabel metal2 s 197624 0 197680 400 6 la_data_in[81]
port 159 nsew signal input
rlabel metal2 s 199304 0 199360 400 6 la_data_in[82]
port 160 nsew signal input
rlabel metal2 s 200984 0 201040 400 6 la_data_in[83]
port 161 nsew signal input
rlabel metal2 s 202664 0 202720 400 6 la_data_in[84]
port 162 nsew signal input
rlabel metal2 s 204344 0 204400 400 6 la_data_in[85]
port 163 nsew signal input
rlabel metal2 s 206024 0 206080 400 6 la_data_in[86]
port 164 nsew signal input
rlabel metal2 s 207704 0 207760 400 6 la_data_in[87]
port 165 nsew signal input
rlabel metal2 s 209384 0 209440 400 6 la_data_in[88]
port 166 nsew signal input
rlabel metal2 s 211064 0 211120 400 6 la_data_in[89]
port 167 nsew signal input
rlabel metal2 s 74984 0 75040 400 6 la_data_in[8]
port 168 nsew signal input
rlabel metal2 s 212744 0 212800 400 6 la_data_in[90]
port 169 nsew signal input
rlabel metal2 s 214424 0 214480 400 6 la_data_in[91]
port 170 nsew signal input
rlabel metal2 s 216104 0 216160 400 6 la_data_in[92]
port 171 nsew signal input
rlabel metal2 s 217784 0 217840 400 6 la_data_in[93]
port 172 nsew signal input
rlabel metal2 s 219464 0 219520 400 6 la_data_in[94]
port 173 nsew signal input
rlabel metal2 s 221144 0 221200 400 6 la_data_in[95]
port 174 nsew signal input
rlabel metal2 s 222824 0 222880 400 6 la_data_in[96]
port 175 nsew signal input
rlabel metal2 s 224504 0 224560 400 6 la_data_in[97]
port 176 nsew signal input
rlabel metal2 s 226184 0 226240 400 6 la_data_in[98]
port 177 nsew signal input
rlabel metal2 s 227864 0 227920 400 6 la_data_in[99]
port 178 nsew signal input
rlabel metal2 s 76664 0 76720 400 6 la_data_in[9]
port 179 nsew signal input
rlabel metal2 s 62104 0 62160 400 6 la_data_out[0]
port 180 nsew signal output
rlabel metal2 s 230104 0 230160 400 6 la_data_out[100]
port 181 nsew signal output
rlabel metal2 s 231784 0 231840 400 6 la_data_out[101]
port 182 nsew signal output
rlabel metal2 s 233464 0 233520 400 6 la_data_out[102]
port 183 nsew signal output
rlabel metal2 s 235144 0 235200 400 6 la_data_out[103]
port 184 nsew signal output
rlabel metal2 s 236824 0 236880 400 6 la_data_out[104]
port 185 nsew signal output
rlabel metal2 s 238504 0 238560 400 6 la_data_out[105]
port 186 nsew signal output
rlabel metal2 s 240184 0 240240 400 6 la_data_out[106]
port 187 nsew signal output
rlabel metal2 s 241864 0 241920 400 6 la_data_out[107]
port 188 nsew signal output
rlabel metal2 s 243544 0 243600 400 6 la_data_out[108]
port 189 nsew signal output
rlabel metal2 s 245224 0 245280 400 6 la_data_out[109]
port 190 nsew signal output
rlabel metal2 s 78904 0 78960 400 6 la_data_out[10]
port 191 nsew signal output
rlabel metal2 s 246904 0 246960 400 6 la_data_out[110]
port 192 nsew signal output
rlabel metal2 s 248584 0 248640 400 6 la_data_out[111]
port 193 nsew signal output
rlabel metal2 s 250264 0 250320 400 6 la_data_out[112]
port 194 nsew signal output
rlabel metal2 s 251944 0 252000 400 6 la_data_out[113]
port 195 nsew signal output
rlabel metal2 s 253624 0 253680 400 6 la_data_out[114]
port 196 nsew signal output
rlabel metal2 s 255304 0 255360 400 6 la_data_out[115]
port 197 nsew signal output
rlabel metal2 s 256984 0 257040 400 6 la_data_out[116]
port 198 nsew signal output
rlabel metal2 s 258664 0 258720 400 6 la_data_out[117]
port 199 nsew signal output
rlabel metal2 s 260344 0 260400 400 6 la_data_out[118]
port 200 nsew signal output
rlabel metal2 s 262024 0 262080 400 6 la_data_out[119]
port 201 nsew signal output
rlabel metal2 s 80584 0 80640 400 6 la_data_out[11]
port 202 nsew signal output
rlabel metal2 s 263704 0 263760 400 6 la_data_out[120]
port 203 nsew signal output
rlabel metal2 s 265384 0 265440 400 6 la_data_out[121]
port 204 nsew signal output
rlabel metal2 s 267064 0 267120 400 6 la_data_out[122]
port 205 nsew signal output
rlabel metal2 s 268744 0 268800 400 6 la_data_out[123]
port 206 nsew signal output
rlabel metal2 s 270424 0 270480 400 6 la_data_out[124]
port 207 nsew signal output
rlabel metal2 s 272104 0 272160 400 6 la_data_out[125]
port 208 nsew signal output
rlabel metal2 s 273784 0 273840 400 6 la_data_out[126]
port 209 nsew signal output
rlabel metal2 s 275464 0 275520 400 6 la_data_out[127]
port 210 nsew signal output
rlabel metal2 s 82264 0 82320 400 6 la_data_out[12]
port 211 nsew signal output
rlabel metal2 s 83944 0 84000 400 6 la_data_out[13]
port 212 nsew signal output
rlabel metal2 s 85624 0 85680 400 6 la_data_out[14]
port 213 nsew signal output
rlabel metal2 s 87304 0 87360 400 6 la_data_out[15]
port 214 nsew signal output
rlabel metal2 s 88984 0 89040 400 6 la_data_out[16]
port 215 nsew signal output
rlabel metal2 s 90664 0 90720 400 6 la_data_out[17]
port 216 nsew signal output
rlabel metal2 s 92344 0 92400 400 6 la_data_out[18]
port 217 nsew signal output
rlabel metal2 s 94024 0 94080 400 6 la_data_out[19]
port 218 nsew signal output
rlabel metal2 s 63784 0 63840 400 6 la_data_out[1]
port 219 nsew signal output
rlabel metal2 s 95704 0 95760 400 6 la_data_out[20]
port 220 nsew signal output
rlabel metal2 s 97384 0 97440 400 6 la_data_out[21]
port 221 nsew signal output
rlabel metal2 s 99064 0 99120 400 6 la_data_out[22]
port 222 nsew signal output
rlabel metal2 s 100744 0 100800 400 6 la_data_out[23]
port 223 nsew signal output
rlabel metal2 s 102424 0 102480 400 6 la_data_out[24]
port 224 nsew signal output
rlabel metal2 s 104104 0 104160 400 6 la_data_out[25]
port 225 nsew signal output
rlabel metal2 s 105784 0 105840 400 6 la_data_out[26]
port 226 nsew signal output
rlabel metal2 s 107464 0 107520 400 6 la_data_out[27]
port 227 nsew signal output
rlabel metal2 s 109144 0 109200 400 6 la_data_out[28]
port 228 nsew signal output
rlabel metal2 s 110824 0 110880 400 6 la_data_out[29]
port 229 nsew signal output
rlabel metal2 s 65464 0 65520 400 6 la_data_out[2]
port 230 nsew signal output
rlabel metal2 s 112504 0 112560 400 6 la_data_out[30]
port 231 nsew signal output
rlabel metal2 s 114184 0 114240 400 6 la_data_out[31]
port 232 nsew signal output
rlabel metal2 s 115864 0 115920 400 6 la_data_out[32]
port 233 nsew signal output
rlabel metal2 s 117544 0 117600 400 6 la_data_out[33]
port 234 nsew signal output
rlabel metal2 s 119224 0 119280 400 6 la_data_out[34]
port 235 nsew signal output
rlabel metal2 s 120904 0 120960 400 6 la_data_out[35]
port 236 nsew signal output
rlabel metal2 s 122584 0 122640 400 6 la_data_out[36]
port 237 nsew signal output
rlabel metal2 s 124264 0 124320 400 6 la_data_out[37]
port 238 nsew signal output
rlabel metal2 s 125944 0 126000 400 6 la_data_out[38]
port 239 nsew signal output
rlabel metal2 s 127624 0 127680 400 6 la_data_out[39]
port 240 nsew signal output
rlabel metal2 s 67144 0 67200 400 6 la_data_out[3]
port 241 nsew signal output
rlabel metal2 s 129304 0 129360 400 6 la_data_out[40]
port 242 nsew signal output
rlabel metal2 s 130984 0 131040 400 6 la_data_out[41]
port 243 nsew signal output
rlabel metal2 s 132664 0 132720 400 6 la_data_out[42]
port 244 nsew signal output
rlabel metal2 s 134344 0 134400 400 6 la_data_out[43]
port 245 nsew signal output
rlabel metal2 s 136024 0 136080 400 6 la_data_out[44]
port 246 nsew signal output
rlabel metal2 s 137704 0 137760 400 6 la_data_out[45]
port 247 nsew signal output
rlabel metal2 s 139384 0 139440 400 6 la_data_out[46]
port 248 nsew signal output
rlabel metal2 s 141064 0 141120 400 6 la_data_out[47]
port 249 nsew signal output
rlabel metal2 s 142744 0 142800 400 6 la_data_out[48]
port 250 nsew signal output
rlabel metal2 s 144424 0 144480 400 6 la_data_out[49]
port 251 nsew signal output
rlabel metal2 s 68824 0 68880 400 6 la_data_out[4]
port 252 nsew signal output
rlabel metal2 s 146104 0 146160 400 6 la_data_out[50]
port 253 nsew signal output
rlabel metal2 s 147784 0 147840 400 6 la_data_out[51]
port 254 nsew signal output
rlabel metal2 s 149464 0 149520 400 6 la_data_out[52]
port 255 nsew signal output
rlabel metal2 s 151144 0 151200 400 6 la_data_out[53]
port 256 nsew signal output
rlabel metal2 s 152824 0 152880 400 6 la_data_out[54]
port 257 nsew signal output
rlabel metal2 s 154504 0 154560 400 6 la_data_out[55]
port 258 nsew signal output
rlabel metal2 s 156184 0 156240 400 6 la_data_out[56]
port 259 nsew signal output
rlabel metal2 s 157864 0 157920 400 6 la_data_out[57]
port 260 nsew signal output
rlabel metal2 s 159544 0 159600 400 6 la_data_out[58]
port 261 nsew signal output
rlabel metal2 s 161224 0 161280 400 6 la_data_out[59]
port 262 nsew signal output
rlabel metal2 s 70504 0 70560 400 6 la_data_out[5]
port 263 nsew signal output
rlabel metal2 s 162904 0 162960 400 6 la_data_out[60]
port 264 nsew signal output
rlabel metal2 s 164584 0 164640 400 6 la_data_out[61]
port 265 nsew signal output
rlabel metal2 s 166264 0 166320 400 6 la_data_out[62]
port 266 nsew signal output
rlabel metal2 s 167944 0 168000 400 6 la_data_out[63]
port 267 nsew signal output
rlabel metal2 s 169624 0 169680 400 6 la_data_out[64]
port 268 nsew signal output
rlabel metal2 s 171304 0 171360 400 6 la_data_out[65]
port 269 nsew signal output
rlabel metal2 s 172984 0 173040 400 6 la_data_out[66]
port 270 nsew signal output
rlabel metal2 s 174664 0 174720 400 6 la_data_out[67]
port 271 nsew signal output
rlabel metal2 s 176344 0 176400 400 6 la_data_out[68]
port 272 nsew signal output
rlabel metal2 s 178024 0 178080 400 6 la_data_out[69]
port 273 nsew signal output
rlabel metal2 s 72184 0 72240 400 6 la_data_out[6]
port 274 nsew signal output
rlabel metal2 s 179704 0 179760 400 6 la_data_out[70]
port 275 nsew signal output
rlabel metal2 s 181384 0 181440 400 6 la_data_out[71]
port 276 nsew signal output
rlabel metal2 s 183064 0 183120 400 6 la_data_out[72]
port 277 nsew signal output
rlabel metal2 s 184744 0 184800 400 6 la_data_out[73]
port 278 nsew signal output
rlabel metal2 s 186424 0 186480 400 6 la_data_out[74]
port 279 nsew signal output
rlabel metal2 s 188104 0 188160 400 6 la_data_out[75]
port 280 nsew signal output
rlabel metal2 s 189784 0 189840 400 6 la_data_out[76]
port 281 nsew signal output
rlabel metal2 s 191464 0 191520 400 6 la_data_out[77]
port 282 nsew signal output
rlabel metal2 s 193144 0 193200 400 6 la_data_out[78]
port 283 nsew signal output
rlabel metal2 s 194824 0 194880 400 6 la_data_out[79]
port 284 nsew signal output
rlabel metal2 s 73864 0 73920 400 6 la_data_out[7]
port 285 nsew signal output
rlabel metal2 s 196504 0 196560 400 6 la_data_out[80]
port 286 nsew signal output
rlabel metal2 s 198184 0 198240 400 6 la_data_out[81]
port 287 nsew signal output
rlabel metal2 s 199864 0 199920 400 6 la_data_out[82]
port 288 nsew signal output
rlabel metal2 s 201544 0 201600 400 6 la_data_out[83]
port 289 nsew signal output
rlabel metal2 s 203224 0 203280 400 6 la_data_out[84]
port 290 nsew signal output
rlabel metal2 s 204904 0 204960 400 6 la_data_out[85]
port 291 nsew signal output
rlabel metal2 s 206584 0 206640 400 6 la_data_out[86]
port 292 nsew signal output
rlabel metal2 s 208264 0 208320 400 6 la_data_out[87]
port 293 nsew signal output
rlabel metal2 s 209944 0 210000 400 6 la_data_out[88]
port 294 nsew signal output
rlabel metal2 s 211624 0 211680 400 6 la_data_out[89]
port 295 nsew signal output
rlabel metal2 s 75544 0 75600 400 6 la_data_out[8]
port 296 nsew signal output
rlabel metal2 s 213304 0 213360 400 6 la_data_out[90]
port 297 nsew signal output
rlabel metal2 s 214984 0 215040 400 6 la_data_out[91]
port 298 nsew signal output
rlabel metal2 s 216664 0 216720 400 6 la_data_out[92]
port 299 nsew signal output
rlabel metal2 s 218344 0 218400 400 6 la_data_out[93]
port 300 nsew signal output
rlabel metal2 s 220024 0 220080 400 6 la_data_out[94]
port 301 nsew signal output
rlabel metal2 s 221704 0 221760 400 6 la_data_out[95]
port 302 nsew signal output
rlabel metal2 s 223384 0 223440 400 6 la_data_out[96]
port 303 nsew signal output
rlabel metal2 s 225064 0 225120 400 6 la_data_out[97]
port 304 nsew signal output
rlabel metal2 s 226744 0 226800 400 6 la_data_out[98]
port 305 nsew signal output
rlabel metal2 s 228424 0 228480 400 6 la_data_out[99]
port 306 nsew signal output
rlabel metal2 s 77224 0 77280 400 6 la_data_out[9]
port 307 nsew signal output
rlabel metal2 s 62664 0 62720 400 6 la_oenb[0]
port 308 nsew signal input
rlabel metal2 s 230664 0 230720 400 6 la_oenb[100]
port 309 nsew signal input
rlabel metal2 s 232344 0 232400 400 6 la_oenb[101]
port 310 nsew signal input
rlabel metal2 s 234024 0 234080 400 6 la_oenb[102]
port 311 nsew signal input
rlabel metal2 s 235704 0 235760 400 6 la_oenb[103]
port 312 nsew signal input
rlabel metal2 s 237384 0 237440 400 6 la_oenb[104]
port 313 nsew signal input
rlabel metal2 s 239064 0 239120 400 6 la_oenb[105]
port 314 nsew signal input
rlabel metal2 s 240744 0 240800 400 6 la_oenb[106]
port 315 nsew signal input
rlabel metal2 s 242424 0 242480 400 6 la_oenb[107]
port 316 nsew signal input
rlabel metal2 s 244104 0 244160 400 6 la_oenb[108]
port 317 nsew signal input
rlabel metal2 s 245784 0 245840 400 6 la_oenb[109]
port 318 nsew signal input
rlabel metal2 s 79464 0 79520 400 6 la_oenb[10]
port 319 nsew signal input
rlabel metal2 s 247464 0 247520 400 6 la_oenb[110]
port 320 nsew signal input
rlabel metal2 s 249144 0 249200 400 6 la_oenb[111]
port 321 nsew signal input
rlabel metal2 s 250824 0 250880 400 6 la_oenb[112]
port 322 nsew signal input
rlabel metal2 s 252504 0 252560 400 6 la_oenb[113]
port 323 nsew signal input
rlabel metal2 s 254184 0 254240 400 6 la_oenb[114]
port 324 nsew signal input
rlabel metal2 s 255864 0 255920 400 6 la_oenb[115]
port 325 nsew signal input
rlabel metal2 s 257544 0 257600 400 6 la_oenb[116]
port 326 nsew signal input
rlabel metal2 s 259224 0 259280 400 6 la_oenb[117]
port 327 nsew signal input
rlabel metal2 s 260904 0 260960 400 6 la_oenb[118]
port 328 nsew signal input
rlabel metal2 s 262584 0 262640 400 6 la_oenb[119]
port 329 nsew signal input
rlabel metal2 s 81144 0 81200 400 6 la_oenb[11]
port 330 nsew signal input
rlabel metal2 s 264264 0 264320 400 6 la_oenb[120]
port 331 nsew signal input
rlabel metal2 s 265944 0 266000 400 6 la_oenb[121]
port 332 nsew signal input
rlabel metal2 s 267624 0 267680 400 6 la_oenb[122]
port 333 nsew signal input
rlabel metal2 s 269304 0 269360 400 6 la_oenb[123]
port 334 nsew signal input
rlabel metal2 s 270984 0 271040 400 6 la_oenb[124]
port 335 nsew signal input
rlabel metal2 s 272664 0 272720 400 6 la_oenb[125]
port 336 nsew signal input
rlabel metal2 s 274344 0 274400 400 6 la_oenb[126]
port 337 nsew signal input
rlabel metal2 s 276024 0 276080 400 6 la_oenb[127]
port 338 nsew signal input
rlabel metal2 s 82824 0 82880 400 6 la_oenb[12]
port 339 nsew signal input
rlabel metal2 s 84504 0 84560 400 6 la_oenb[13]
port 340 nsew signal input
rlabel metal2 s 86184 0 86240 400 6 la_oenb[14]
port 341 nsew signal input
rlabel metal2 s 87864 0 87920 400 6 la_oenb[15]
port 342 nsew signal input
rlabel metal2 s 89544 0 89600 400 6 la_oenb[16]
port 343 nsew signal input
rlabel metal2 s 91224 0 91280 400 6 la_oenb[17]
port 344 nsew signal input
rlabel metal2 s 92904 0 92960 400 6 la_oenb[18]
port 345 nsew signal input
rlabel metal2 s 94584 0 94640 400 6 la_oenb[19]
port 346 nsew signal input
rlabel metal2 s 64344 0 64400 400 6 la_oenb[1]
port 347 nsew signal input
rlabel metal2 s 96264 0 96320 400 6 la_oenb[20]
port 348 nsew signal input
rlabel metal2 s 97944 0 98000 400 6 la_oenb[21]
port 349 nsew signal input
rlabel metal2 s 99624 0 99680 400 6 la_oenb[22]
port 350 nsew signal input
rlabel metal2 s 101304 0 101360 400 6 la_oenb[23]
port 351 nsew signal input
rlabel metal2 s 102984 0 103040 400 6 la_oenb[24]
port 352 nsew signal input
rlabel metal2 s 104664 0 104720 400 6 la_oenb[25]
port 353 nsew signal input
rlabel metal2 s 106344 0 106400 400 6 la_oenb[26]
port 354 nsew signal input
rlabel metal2 s 108024 0 108080 400 6 la_oenb[27]
port 355 nsew signal input
rlabel metal2 s 109704 0 109760 400 6 la_oenb[28]
port 356 nsew signal input
rlabel metal2 s 111384 0 111440 400 6 la_oenb[29]
port 357 nsew signal input
rlabel metal2 s 66024 0 66080 400 6 la_oenb[2]
port 358 nsew signal input
rlabel metal2 s 113064 0 113120 400 6 la_oenb[30]
port 359 nsew signal input
rlabel metal2 s 114744 0 114800 400 6 la_oenb[31]
port 360 nsew signal input
rlabel metal2 s 116424 0 116480 400 6 la_oenb[32]
port 361 nsew signal input
rlabel metal2 s 118104 0 118160 400 6 la_oenb[33]
port 362 nsew signal input
rlabel metal2 s 119784 0 119840 400 6 la_oenb[34]
port 363 nsew signal input
rlabel metal2 s 121464 0 121520 400 6 la_oenb[35]
port 364 nsew signal input
rlabel metal2 s 123144 0 123200 400 6 la_oenb[36]
port 365 nsew signal input
rlabel metal2 s 124824 0 124880 400 6 la_oenb[37]
port 366 nsew signal input
rlabel metal2 s 126504 0 126560 400 6 la_oenb[38]
port 367 nsew signal input
rlabel metal2 s 128184 0 128240 400 6 la_oenb[39]
port 368 nsew signal input
rlabel metal2 s 67704 0 67760 400 6 la_oenb[3]
port 369 nsew signal input
rlabel metal2 s 129864 0 129920 400 6 la_oenb[40]
port 370 nsew signal input
rlabel metal2 s 131544 0 131600 400 6 la_oenb[41]
port 371 nsew signal input
rlabel metal2 s 133224 0 133280 400 6 la_oenb[42]
port 372 nsew signal input
rlabel metal2 s 134904 0 134960 400 6 la_oenb[43]
port 373 nsew signal input
rlabel metal2 s 136584 0 136640 400 6 la_oenb[44]
port 374 nsew signal input
rlabel metal2 s 138264 0 138320 400 6 la_oenb[45]
port 375 nsew signal input
rlabel metal2 s 139944 0 140000 400 6 la_oenb[46]
port 376 nsew signal input
rlabel metal2 s 141624 0 141680 400 6 la_oenb[47]
port 377 nsew signal input
rlabel metal2 s 143304 0 143360 400 6 la_oenb[48]
port 378 nsew signal input
rlabel metal2 s 144984 0 145040 400 6 la_oenb[49]
port 379 nsew signal input
rlabel metal2 s 69384 0 69440 400 6 la_oenb[4]
port 380 nsew signal input
rlabel metal2 s 146664 0 146720 400 6 la_oenb[50]
port 381 nsew signal input
rlabel metal2 s 148344 0 148400 400 6 la_oenb[51]
port 382 nsew signal input
rlabel metal2 s 150024 0 150080 400 6 la_oenb[52]
port 383 nsew signal input
rlabel metal2 s 151704 0 151760 400 6 la_oenb[53]
port 384 nsew signal input
rlabel metal2 s 153384 0 153440 400 6 la_oenb[54]
port 385 nsew signal input
rlabel metal2 s 155064 0 155120 400 6 la_oenb[55]
port 386 nsew signal input
rlabel metal2 s 156744 0 156800 400 6 la_oenb[56]
port 387 nsew signal input
rlabel metal2 s 158424 0 158480 400 6 la_oenb[57]
port 388 nsew signal input
rlabel metal2 s 160104 0 160160 400 6 la_oenb[58]
port 389 nsew signal input
rlabel metal2 s 161784 0 161840 400 6 la_oenb[59]
port 390 nsew signal input
rlabel metal2 s 71064 0 71120 400 6 la_oenb[5]
port 391 nsew signal input
rlabel metal2 s 163464 0 163520 400 6 la_oenb[60]
port 392 nsew signal input
rlabel metal2 s 165144 0 165200 400 6 la_oenb[61]
port 393 nsew signal input
rlabel metal2 s 166824 0 166880 400 6 la_oenb[62]
port 394 nsew signal input
rlabel metal2 s 168504 0 168560 400 6 la_oenb[63]
port 395 nsew signal input
rlabel metal2 s 170184 0 170240 400 6 la_oenb[64]
port 396 nsew signal input
rlabel metal2 s 171864 0 171920 400 6 la_oenb[65]
port 397 nsew signal input
rlabel metal2 s 173544 0 173600 400 6 la_oenb[66]
port 398 nsew signal input
rlabel metal2 s 175224 0 175280 400 6 la_oenb[67]
port 399 nsew signal input
rlabel metal2 s 176904 0 176960 400 6 la_oenb[68]
port 400 nsew signal input
rlabel metal2 s 178584 0 178640 400 6 la_oenb[69]
port 401 nsew signal input
rlabel metal2 s 72744 0 72800 400 6 la_oenb[6]
port 402 nsew signal input
rlabel metal2 s 180264 0 180320 400 6 la_oenb[70]
port 403 nsew signal input
rlabel metal2 s 181944 0 182000 400 6 la_oenb[71]
port 404 nsew signal input
rlabel metal2 s 183624 0 183680 400 6 la_oenb[72]
port 405 nsew signal input
rlabel metal2 s 185304 0 185360 400 6 la_oenb[73]
port 406 nsew signal input
rlabel metal2 s 186984 0 187040 400 6 la_oenb[74]
port 407 nsew signal input
rlabel metal2 s 188664 0 188720 400 6 la_oenb[75]
port 408 nsew signal input
rlabel metal2 s 190344 0 190400 400 6 la_oenb[76]
port 409 nsew signal input
rlabel metal2 s 192024 0 192080 400 6 la_oenb[77]
port 410 nsew signal input
rlabel metal2 s 193704 0 193760 400 6 la_oenb[78]
port 411 nsew signal input
rlabel metal2 s 195384 0 195440 400 6 la_oenb[79]
port 412 nsew signal input
rlabel metal2 s 74424 0 74480 400 6 la_oenb[7]
port 413 nsew signal input
rlabel metal2 s 197064 0 197120 400 6 la_oenb[80]
port 414 nsew signal input
rlabel metal2 s 198744 0 198800 400 6 la_oenb[81]
port 415 nsew signal input
rlabel metal2 s 200424 0 200480 400 6 la_oenb[82]
port 416 nsew signal input
rlabel metal2 s 202104 0 202160 400 6 la_oenb[83]
port 417 nsew signal input
rlabel metal2 s 203784 0 203840 400 6 la_oenb[84]
port 418 nsew signal input
rlabel metal2 s 205464 0 205520 400 6 la_oenb[85]
port 419 nsew signal input
rlabel metal2 s 207144 0 207200 400 6 la_oenb[86]
port 420 nsew signal input
rlabel metal2 s 208824 0 208880 400 6 la_oenb[87]
port 421 nsew signal input
rlabel metal2 s 210504 0 210560 400 6 la_oenb[88]
port 422 nsew signal input
rlabel metal2 s 212184 0 212240 400 6 la_oenb[89]
port 423 nsew signal input
rlabel metal2 s 76104 0 76160 400 6 la_oenb[8]
port 424 nsew signal input
rlabel metal2 s 213864 0 213920 400 6 la_oenb[90]
port 425 nsew signal input
rlabel metal2 s 215544 0 215600 400 6 la_oenb[91]
port 426 nsew signal input
rlabel metal2 s 217224 0 217280 400 6 la_oenb[92]
port 427 nsew signal input
rlabel metal2 s 218904 0 218960 400 6 la_oenb[93]
port 428 nsew signal input
rlabel metal2 s 220584 0 220640 400 6 la_oenb[94]
port 429 nsew signal input
rlabel metal2 s 222264 0 222320 400 6 la_oenb[95]
port 430 nsew signal input
rlabel metal2 s 223944 0 224000 400 6 la_oenb[96]
port 431 nsew signal input
rlabel metal2 s 225624 0 225680 400 6 la_oenb[97]
port 432 nsew signal input
rlabel metal2 s 227304 0 227360 400 6 la_oenb[98]
port 433 nsew signal input
rlabel metal2 s 228984 0 229040 400 6 la_oenb[99]
port 434 nsew signal input
rlabel metal2 s 77784 0 77840 400 6 la_oenb[9]
port 435 nsew signal input
rlabel metal4 s 2224 1538 2384 174078 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 174078 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 174078 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 174078 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 174078 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 174078 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 174078 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 174078 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 174078 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 174078 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 174078 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 174078 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 174078 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 174078 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 174078 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 174078 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 174078 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 263344 1538 263504 174078 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 278704 1538 278864 174078 6 vccd1
port 436 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 174078 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 174078 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 174078 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 174078 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 174078 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 174078 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 174078 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 174078 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 174078 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 174078 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 174078 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 174078 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 174078 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 174078 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 174078 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 174078 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 255664 1538 255824 174078 6 vssd1
port 437 nsew ground bidirectional
rlabel metal4 s 271024 1538 271184 174078 6 vssd1
port 437 nsew ground bidirectional
rlabel metal2 s 2184 0 2240 400 6 wb_clk_i
port 438 nsew signal input
rlabel metal2 s 2744 0 2800 400 6 wb_rst_i
port 439 nsew signal input
rlabel metal2 s 3304 0 3360 400 6 wbs_ack_o
port 440 nsew signal output
rlabel metal2 s 5544 0 5600 400 6 wbs_adr_i[0]
port 441 nsew signal input
rlabel metal2 s 24584 0 24640 400 6 wbs_adr_i[10]
port 442 nsew signal input
rlabel metal2 s 26264 0 26320 400 6 wbs_adr_i[11]
port 443 nsew signal input
rlabel metal2 s 27944 0 28000 400 6 wbs_adr_i[12]
port 444 nsew signal input
rlabel metal2 s 29624 0 29680 400 6 wbs_adr_i[13]
port 445 nsew signal input
rlabel metal2 s 31304 0 31360 400 6 wbs_adr_i[14]
port 446 nsew signal input
rlabel metal2 s 32984 0 33040 400 6 wbs_adr_i[15]
port 447 nsew signal input
rlabel metal2 s 34664 0 34720 400 6 wbs_adr_i[16]
port 448 nsew signal input
rlabel metal2 s 36344 0 36400 400 6 wbs_adr_i[17]
port 449 nsew signal input
rlabel metal2 s 38024 0 38080 400 6 wbs_adr_i[18]
port 450 nsew signal input
rlabel metal2 s 39704 0 39760 400 6 wbs_adr_i[19]
port 451 nsew signal input
rlabel metal2 s 7784 0 7840 400 6 wbs_adr_i[1]
port 452 nsew signal input
rlabel metal2 s 41384 0 41440 400 6 wbs_adr_i[20]
port 453 nsew signal input
rlabel metal2 s 43064 0 43120 400 6 wbs_adr_i[21]
port 454 nsew signal input
rlabel metal2 s 44744 0 44800 400 6 wbs_adr_i[22]
port 455 nsew signal input
rlabel metal2 s 46424 0 46480 400 6 wbs_adr_i[23]
port 456 nsew signal input
rlabel metal2 s 48104 0 48160 400 6 wbs_adr_i[24]
port 457 nsew signal input
rlabel metal2 s 49784 0 49840 400 6 wbs_adr_i[25]
port 458 nsew signal input
rlabel metal2 s 51464 0 51520 400 6 wbs_adr_i[26]
port 459 nsew signal input
rlabel metal2 s 53144 0 53200 400 6 wbs_adr_i[27]
port 460 nsew signal input
rlabel metal2 s 54824 0 54880 400 6 wbs_adr_i[28]
port 461 nsew signal input
rlabel metal2 s 56504 0 56560 400 6 wbs_adr_i[29]
port 462 nsew signal input
rlabel metal2 s 10024 0 10080 400 6 wbs_adr_i[2]
port 463 nsew signal input
rlabel metal2 s 58184 0 58240 400 6 wbs_adr_i[30]
port 464 nsew signal input
rlabel metal2 s 59864 0 59920 400 6 wbs_adr_i[31]
port 465 nsew signal input
rlabel metal2 s 12264 0 12320 400 6 wbs_adr_i[3]
port 466 nsew signal input
rlabel metal2 s 14504 0 14560 400 6 wbs_adr_i[4]
port 467 nsew signal input
rlabel metal2 s 16184 0 16240 400 6 wbs_adr_i[5]
port 468 nsew signal input
rlabel metal2 s 17864 0 17920 400 6 wbs_adr_i[6]
port 469 nsew signal input
rlabel metal2 s 19544 0 19600 400 6 wbs_adr_i[7]
port 470 nsew signal input
rlabel metal2 s 21224 0 21280 400 6 wbs_adr_i[8]
port 471 nsew signal input
rlabel metal2 s 22904 0 22960 400 6 wbs_adr_i[9]
port 472 nsew signal input
rlabel metal2 s 3864 0 3920 400 6 wbs_cyc_i
port 473 nsew signal input
rlabel metal2 s 6104 0 6160 400 6 wbs_dat_i[0]
port 474 nsew signal input
rlabel metal2 s 25144 0 25200 400 6 wbs_dat_i[10]
port 475 nsew signal input
rlabel metal2 s 26824 0 26880 400 6 wbs_dat_i[11]
port 476 nsew signal input
rlabel metal2 s 28504 0 28560 400 6 wbs_dat_i[12]
port 477 nsew signal input
rlabel metal2 s 30184 0 30240 400 6 wbs_dat_i[13]
port 478 nsew signal input
rlabel metal2 s 31864 0 31920 400 6 wbs_dat_i[14]
port 479 nsew signal input
rlabel metal2 s 33544 0 33600 400 6 wbs_dat_i[15]
port 480 nsew signal input
rlabel metal2 s 35224 0 35280 400 6 wbs_dat_i[16]
port 481 nsew signal input
rlabel metal2 s 36904 0 36960 400 6 wbs_dat_i[17]
port 482 nsew signal input
rlabel metal2 s 38584 0 38640 400 6 wbs_dat_i[18]
port 483 nsew signal input
rlabel metal2 s 40264 0 40320 400 6 wbs_dat_i[19]
port 484 nsew signal input
rlabel metal2 s 8344 0 8400 400 6 wbs_dat_i[1]
port 485 nsew signal input
rlabel metal2 s 41944 0 42000 400 6 wbs_dat_i[20]
port 486 nsew signal input
rlabel metal2 s 43624 0 43680 400 6 wbs_dat_i[21]
port 487 nsew signal input
rlabel metal2 s 45304 0 45360 400 6 wbs_dat_i[22]
port 488 nsew signal input
rlabel metal2 s 46984 0 47040 400 6 wbs_dat_i[23]
port 489 nsew signal input
rlabel metal2 s 48664 0 48720 400 6 wbs_dat_i[24]
port 490 nsew signal input
rlabel metal2 s 50344 0 50400 400 6 wbs_dat_i[25]
port 491 nsew signal input
rlabel metal2 s 52024 0 52080 400 6 wbs_dat_i[26]
port 492 nsew signal input
rlabel metal2 s 53704 0 53760 400 6 wbs_dat_i[27]
port 493 nsew signal input
rlabel metal2 s 55384 0 55440 400 6 wbs_dat_i[28]
port 494 nsew signal input
rlabel metal2 s 57064 0 57120 400 6 wbs_dat_i[29]
port 495 nsew signal input
rlabel metal2 s 10584 0 10640 400 6 wbs_dat_i[2]
port 496 nsew signal input
rlabel metal2 s 58744 0 58800 400 6 wbs_dat_i[30]
port 497 nsew signal input
rlabel metal2 s 60424 0 60480 400 6 wbs_dat_i[31]
port 498 nsew signal input
rlabel metal2 s 12824 0 12880 400 6 wbs_dat_i[3]
port 499 nsew signal input
rlabel metal2 s 15064 0 15120 400 6 wbs_dat_i[4]
port 500 nsew signal input
rlabel metal2 s 16744 0 16800 400 6 wbs_dat_i[5]
port 501 nsew signal input
rlabel metal2 s 18424 0 18480 400 6 wbs_dat_i[6]
port 502 nsew signal input
rlabel metal2 s 20104 0 20160 400 6 wbs_dat_i[7]
port 503 nsew signal input
rlabel metal2 s 21784 0 21840 400 6 wbs_dat_i[8]
port 504 nsew signal input
rlabel metal2 s 23464 0 23520 400 6 wbs_dat_i[9]
port 505 nsew signal input
rlabel metal2 s 6664 0 6720 400 6 wbs_dat_o[0]
port 506 nsew signal output
rlabel metal2 s 25704 0 25760 400 6 wbs_dat_o[10]
port 507 nsew signal output
rlabel metal2 s 27384 0 27440 400 6 wbs_dat_o[11]
port 508 nsew signal output
rlabel metal2 s 29064 0 29120 400 6 wbs_dat_o[12]
port 509 nsew signal output
rlabel metal2 s 30744 0 30800 400 6 wbs_dat_o[13]
port 510 nsew signal output
rlabel metal2 s 32424 0 32480 400 6 wbs_dat_o[14]
port 511 nsew signal output
rlabel metal2 s 34104 0 34160 400 6 wbs_dat_o[15]
port 512 nsew signal output
rlabel metal2 s 35784 0 35840 400 6 wbs_dat_o[16]
port 513 nsew signal output
rlabel metal2 s 37464 0 37520 400 6 wbs_dat_o[17]
port 514 nsew signal output
rlabel metal2 s 39144 0 39200 400 6 wbs_dat_o[18]
port 515 nsew signal output
rlabel metal2 s 40824 0 40880 400 6 wbs_dat_o[19]
port 516 nsew signal output
rlabel metal2 s 8904 0 8960 400 6 wbs_dat_o[1]
port 517 nsew signal output
rlabel metal2 s 42504 0 42560 400 6 wbs_dat_o[20]
port 518 nsew signal output
rlabel metal2 s 44184 0 44240 400 6 wbs_dat_o[21]
port 519 nsew signal output
rlabel metal2 s 45864 0 45920 400 6 wbs_dat_o[22]
port 520 nsew signal output
rlabel metal2 s 47544 0 47600 400 6 wbs_dat_o[23]
port 521 nsew signal output
rlabel metal2 s 49224 0 49280 400 6 wbs_dat_o[24]
port 522 nsew signal output
rlabel metal2 s 50904 0 50960 400 6 wbs_dat_o[25]
port 523 nsew signal output
rlabel metal2 s 52584 0 52640 400 6 wbs_dat_o[26]
port 524 nsew signal output
rlabel metal2 s 54264 0 54320 400 6 wbs_dat_o[27]
port 525 nsew signal output
rlabel metal2 s 55944 0 56000 400 6 wbs_dat_o[28]
port 526 nsew signal output
rlabel metal2 s 57624 0 57680 400 6 wbs_dat_o[29]
port 527 nsew signal output
rlabel metal2 s 11144 0 11200 400 6 wbs_dat_o[2]
port 528 nsew signal output
rlabel metal2 s 59304 0 59360 400 6 wbs_dat_o[30]
port 529 nsew signal output
rlabel metal2 s 60984 0 61040 400 6 wbs_dat_o[31]
port 530 nsew signal output
rlabel metal2 s 13384 0 13440 400 6 wbs_dat_o[3]
port 531 nsew signal output
rlabel metal2 s 15624 0 15680 400 6 wbs_dat_o[4]
port 532 nsew signal output
rlabel metal2 s 17304 0 17360 400 6 wbs_dat_o[5]
port 533 nsew signal output
rlabel metal2 s 18984 0 19040 400 6 wbs_dat_o[6]
port 534 nsew signal output
rlabel metal2 s 20664 0 20720 400 6 wbs_dat_o[7]
port 535 nsew signal output
rlabel metal2 s 22344 0 22400 400 6 wbs_dat_o[8]
port 536 nsew signal output
rlabel metal2 s 24024 0 24080 400 6 wbs_dat_o[9]
port 537 nsew signal output
rlabel metal2 s 7224 0 7280 400 6 wbs_sel_i[0]
port 538 nsew signal input
rlabel metal2 s 9464 0 9520 400 6 wbs_sel_i[1]
port 539 nsew signal input
rlabel metal2 s 11704 0 11760 400 6 wbs_sel_i[2]
port 540 nsew signal input
rlabel metal2 s 13944 0 14000 400 6 wbs_sel_i[3]
port 541 nsew signal input
rlabel metal2 s 4424 0 4480 400 6 wbs_stb_i
port 542 nsew signal input
rlabel metal2 s 4984 0 5040 400 6 wbs_we_i
port 543 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 280000 176000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17708586
string GDS_FILE /home/sangamanath/Desktop/ring_counter_caravel/openlane/user_proj_example/runs/23_07_10_15_44/results/signoff/user_proj_example.magic.gds
string GDS_START 297514
<< end >>

