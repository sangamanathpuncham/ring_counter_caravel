module ring_counter (Clock,
    Reset,
    vccd1,
    vssd1,
    Count_out,
    io_oeb);
 input Clock;
 input Reset;
 input vccd1;
 input vssd1;
 output [3:0] Count_out;
 output [3:0] io_oeb;

 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire clknet_0_Clock;
 wire clknet_1_0__leaf_Clock;
 wire clknet_1_1__leaf_Clock;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;

 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_19 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_187 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_191 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_242 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_160 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_164 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_166 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_214 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_246 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_196 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_202 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_220 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_231 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_160 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_195 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_201 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_294 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_298 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_305 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_23 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_31 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_7 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_104 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_107 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_139 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_142 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_174 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_177 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_18 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_197 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_205 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_209 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_23 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_244 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_282 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_31 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_317 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_325 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_69 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_72 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_321 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_329 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_286 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_318 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_326 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_330 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 (.VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_110 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_111 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_112 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_113 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_114 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_115 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_116 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_117 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_118 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_119 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_120 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_121 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_122 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_123 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_124 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_125 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_126 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_127 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_128 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_129 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_130 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_131 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_132 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_133 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_134 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_135 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_136 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_138 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_139 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_140 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_142 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_143 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_145 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_146 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_147 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_148 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_149 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_150 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_151 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_152 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_153 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_154 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_155 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_156 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_157 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_158 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_159 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_160 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_161 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_162 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_163 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_164 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_165 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_166 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_167 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_168 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_169 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_170 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_171 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_173 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_174 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_175 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_177 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_178 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_180 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_181 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_182 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_183 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_184 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_185 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_186 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_187 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _04_ (.I(net1),
    .ZN(_00_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05_ (.I(net1),
    .ZN(_01_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06_ (.I(net1),
    .ZN(_02_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07_ (.I(net1),
    .ZN(_03_),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _08_ (.D(net5),
    .SETN(_00_),
    .CLK(clknet_1_0__leaf_Clock),
    .Q(net2),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _09_ (.D(net2),
    .RN(_01_),
    .CLK(clknet_1_0__leaf_Clock),
    .Q(net3),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _10_ (.D(net3),
    .RN(_02_),
    .CLK(clknet_1_1__leaf_Clock),
    .Q(net4),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _11_ (.D(net4),
    .RN(_03_),
    .CLK(clknet_1_1__leaf_Clock),
    .Q(net5),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_Clock (.I(Clock),
    .Z(clknet_0_Clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_Clock (.I(clknet_0_Clock),
    .Z(clknet_1_0__leaf_Clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_Clock (.I(clknet_0_Clock),
    .Z(clknet_1_1__leaf_Clock),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1 (.I(Reset),
    .Z(net1),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output2 (.I(net2),
    .Z(Count_out[0]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output3 (.I(net3),
    .Z(Count_out[1]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output4 (.I(net4),
    .Z(Count_out[2]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output5 (.I(net5),
    .Z(Count_out[3]),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel ring_counter_6 (.ZN(net6),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel ring_counter_7 (.ZN(net7),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel ring_counter_8 (.ZN(net8),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel ring_counter_9 (.ZN(net9),
    .VDD(vccd1),
    .VNW(vccd1),
    .VPW(vssd1),
    .VSS(vssd1));
 assign io_oeb[0] = net6;
 assign io_oeb[1] = net7;
 assign io_oeb[2] = net8;
 assign io_oeb[3] = net9;
endmodule
